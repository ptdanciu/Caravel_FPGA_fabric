(* blackbox *) module rram_28(
	input WL,
    input [0:27] BL,
    output [0:27] Q
);
endmodule
