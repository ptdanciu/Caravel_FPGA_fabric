module test_lut_inst (clk,
    data_in,
    enable,
    reset,
    set,
    bl_address,
    gfpga_pad_GPIO_PAD,
    wl_address);
 input clk;
 input data_in;
 input enable;
 input reset;
 input set;
 input [4:0] bl_address;
 inout [31:0] gfpga_pad_GPIO_PAD;
 input [4:0] wl_address;

 wire VDD;
 wire VSS;
 wire \Q27[10] ;
 wire \Q27[11] ;
 wire \Q27[12] ;
 wire \Q27[13] ;
 wire \Q27[14] ;
 wire \Q27[15] ;
 wire \Q27[16] ;
 wire \Q27[17] ;
 wire \Q27[18] ;
 wire \Q27[19] ;
 wire \Q27[20] ;
 wire \Q27[21] ;
 wire \Q27[22] ;
 wire \Q27[23] ;
 wire \Q27[24] ;
 wire \Q27[25] ;
 wire \Q27[26] ;
 wire \Q27[27] ;
 wire \Q27[28] ;
 wire \Q27[7] ;
 wire \Q27[8] ;
 wire \Q27[9] ;
 wire \Q5[13] ;
 wire \Q5[14] ;
 wire \Q5[15] ;
 wire \Q5[16] ;
 wire \Q5[17] ;
 wire \Q5[18] ;
 wire \Q5[19] ;
 wire \Q5[20] ;
 wire \Q5[21] ;
 wire \Q5[22] ;
 wire \Q5[23] ;
 wire \Q5[24] ;
 wire \Q5[25] ;
 wire \Q5[26] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0588_;
 wire _0589_;
 wire _0592_;
 wire _0593_;
 wire _0595_;
 wire _0598_;
 wire _0599_;
 wire _0601_;
 wire _0602_;
 wire _0604_;
 wire _0605_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire \cbx_1__0_.Q_in[0] ;
 wire \cbx_1__0_.Q_in[10] ;
 wire \cbx_1__0_.Q_in[11] ;
 wire \cbx_1__0_.Q_in[12] ;
 wire \cbx_1__0_.Q_in[13] ;
 wire \cbx_1__0_.Q_in[14] ;
 wire \cbx_1__0_.Q_in[15] ;
 wire \cbx_1__0_.Q_in[16] ;
 wire \cbx_1__0_.Q_in[17] ;
 wire \cbx_1__0_.Q_in[18] ;
 wire \cbx_1__0_.Q_in[19] ;
 wire \cbx_1__0_.Q_in[1] ;
 wire \cbx_1__0_.Q_in[20] ;
 wire \cbx_1__0_.Q_in[21] ;
 wire \cbx_1__0_.Q_in[22] ;
 wire \cbx_1__0_.Q_in[23] ;
 wire \cbx_1__0_.Q_in[24] ;
 wire \cbx_1__0_.Q_in[25] ;
 wire \cbx_1__0_.Q_in[26] ;
 wire \cbx_1__0_.Q_in[27] ;
 wire \cbx_1__0_.Q_in[28] ;
 wire \cbx_1__0_.Q_in[29] ;
 wire \cbx_1__0_.Q_in[2] ;
 wire \cbx_1__0_.Q_in[30] ;
 wire \cbx_1__0_.Q_in[31] ;
 wire \cbx_1__0_.Q_in[32] ;
 wire \cbx_1__0_.Q_in[33] ;
 wire \cbx_1__0_.Q_in[34] ;
 wire \cbx_1__0_.Q_in[35] ;
 wire \cbx_1__0_.Q_in[36] ;
 wire \cbx_1__0_.Q_in[37] ;
 wire \cbx_1__0_.Q_in[38] ;
 wire \cbx_1__0_.Q_in[39] ;
 wire \cbx_1__0_.Q_in[3] ;
 wire \cbx_1__0_.Q_in[40] ;
 wire \cbx_1__0_.Q_in[41] ;
 wire \cbx_1__0_.Q_in[42] ;
 wire \cbx_1__0_.Q_in[43] ;
 wire \cbx_1__0_.Q_in[44] ;
 wire \cbx_1__0_.Q_in[45] ;
 wire \cbx_1__0_.Q_in[46] ;
 wire \cbx_1__0_.Q_in[47] ;
 wire \cbx_1__0_.Q_in[48] ;
 wire \cbx_1__0_.Q_in[49] ;
 wire \cbx_1__0_.Q_in[4] ;
 wire \cbx_1__0_.Q_in[50] ;
 wire \cbx_1__0_.Q_in[51] ;
 wire \cbx_1__0_.Q_in[52] ;
 wire \cbx_1__0_.Q_in[53] ;
 wire \cbx_1__0_.Q_in[54] ;
 wire \cbx_1__0_.Q_in[55] ;
 wire \cbx_1__0_.Q_in[56] ;
 wire \cbx_1__0_.Q_in[57] ;
 wire \cbx_1__0_.Q_in[58] ;
 wire \cbx_1__0_.Q_in[59] ;
 wire \cbx_1__0_.Q_in[5] ;
 wire \cbx_1__0_.Q_in[60] ;
 wire \cbx_1__0_.Q_in[61] ;
 wire \cbx_1__0_.Q_in[62] ;
 wire \cbx_1__0_.Q_in[63] ;
 wire \cbx_1__0_.Q_in[64] ;
 wire \cbx_1__0_.Q_in[65] ;
 wire \cbx_1__0_.Q_in[6] ;
 wire \cbx_1__0_.Q_in[7] ;
 wire \cbx_1__0_.Q_in[8] ;
 wire \cbx_1__0_.Q_in[9] ;
 wire \cbx_1__0_.mux_bottom_ipin_0.INVTX1_4_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.INVTX1_5_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_2.INVTX1_2_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.INVTX1_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.INVTX1_3_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.INVTX1_4_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.INVTX1_5_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.INVTX1_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.INVTX1_3_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.INVTX1_4_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.INVTX1_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.INVTX1_3_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__0_.wl[0] ;
 wire \cbx_1__0_.wl[10] ;
 wire \cbx_1__0_.wl[11] ;
 wire \cbx_1__0_.wl[12] ;
 wire \cbx_1__0_.wl[13] ;
 wire \cbx_1__0_.wl[14] ;
 wire \cbx_1__0_.wl[15] ;
 wire \cbx_1__0_.wl[16] ;
 wire \cbx_1__0_.wl[17] ;
 wire \cbx_1__0_.wl[18] ;
 wire \cbx_1__0_.wl[19] ;
 wire \cbx_1__0_.wl[1] ;
 wire \cbx_1__0_.wl[20] ;
 wire \cbx_1__0_.wl[21] ;
 wire \cbx_1__0_.wl[22] ;
 wire \cbx_1__0_.wl[23] ;
 wire \cbx_1__0_.wl[24] ;
 wire \cbx_1__0_.wl[25] ;
 wire \cbx_1__0_.wl[26] ;
 wire \cbx_1__0_.wl[27] ;
 wire \cbx_1__0_.wl[28] ;
 wire \cbx_1__0_.wl[2] ;
 wire \cbx_1__0_.wl[32] ;
 wire \cbx_1__0_.wl[33] ;
 wire \cbx_1__0_.wl[34] ;
 wire \cbx_1__0_.wl[35] ;
 wire \cbx_1__0_.wl[36] ;
 wire \cbx_1__0_.wl[37] ;
 wire \cbx_1__0_.wl[38] ;
 wire \cbx_1__1_.Q_in[0] ;
 wire \cbx_1__1_.Q_in[10] ;
 wire \cbx_1__1_.Q_in[11] ;
 wire \cbx_1__1_.Q_in[12] ;
 wire \cbx_1__1_.Q_in[13] ;
 wire \cbx_1__1_.Q_in[14] ;
 wire \cbx_1__1_.Q_in[15] ;
 wire \cbx_1__1_.Q_in[16] ;
 wire \cbx_1__1_.Q_in[17] ;
 wire \cbx_1__1_.Q_in[18] ;
 wire \cbx_1__1_.Q_in[19] ;
 wire \cbx_1__1_.Q_in[1] ;
 wire \cbx_1__1_.Q_in[20] ;
 wire \cbx_1__1_.Q_in[21] ;
 wire \cbx_1__1_.Q_in[22] ;
 wire \cbx_1__1_.Q_in[23] ;
 wire \cbx_1__1_.Q_in[24] ;
 wire \cbx_1__1_.Q_in[25] ;
 wire \cbx_1__1_.Q_in[26] ;
 wire \cbx_1__1_.Q_in[27] ;
 wire \cbx_1__1_.Q_in[28] ;
 wire \cbx_1__1_.Q_in[29] ;
 wire \cbx_1__1_.Q_in[2] ;
 wire \cbx_1__1_.Q_in[30] ;
 wire \cbx_1__1_.Q_in[31] ;
 wire \cbx_1__1_.Q_in[32] ;
 wire \cbx_1__1_.Q_in[33] ;
 wire \cbx_1__1_.Q_in[34] ;
 wire \cbx_1__1_.Q_in[35] ;
 wire \cbx_1__1_.Q_in[36] ;
 wire \cbx_1__1_.Q_in[37] ;
 wire \cbx_1__1_.Q_in[38] ;
 wire \cbx_1__1_.Q_in[39] ;
 wire \cbx_1__1_.Q_in[3] ;
 wire \cbx_1__1_.Q_in[40] ;
 wire \cbx_1__1_.Q_in[41] ;
 wire \cbx_1__1_.Q_in[42] ;
 wire \cbx_1__1_.Q_in[43] ;
 wire \cbx_1__1_.Q_in[44] ;
 wire \cbx_1__1_.Q_in[45] ;
 wire \cbx_1__1_.Q_in[46] ;
 wire \cbx_1__1_.Q_in[47] ;
 wire \cbx_1__1_.Q_in[48] ;
 wire \cbx_1__1_.Q_in[49] ;
 wire \cbx_1__1_.Q_in[4] ;
 wire \cbx_1__1_.Q_in[50] ;
 wire \cbx_1__1_.Q_in[51] ;
 wire \cbx_1__1_.Q_in[52] ;
 wire \cbx_1__1_.Q_in[53] ;
 wire \cbx_1__1_.Q_in[54] ;
 wire \cbx_1__1_.Q_in[55] ;
 wire \cbx_1__1_.Q_in[56] ;
 wire \cbx_1__1_.Q_in[57] ;
 wire \cbx_1__1_.Q_in[58] ;
 wire \cbx_1__1_.Q_in[59] ;
 wire \cbx_1__1_.Q_in[5] ;
 wire \cbx_1__1_.Q_in[60] ;
 wire \cbx_1__1_.Q_in[61] ;
 wire \cbx_1__1_.Q_in[62] ;
 wire \cbx_1__1_.Q_in[63] ;
 wire \cbx_1__1_.Q_in[64] ;
 wire \cbx_1__1_.Q_in[65] ;
 wire \cbx_1__1_.Q_in[6] ;
 wire \cbx_1__1_.Q_in[7] ;
 wire \cbx_1__1_.Q_in[8] ;
 wire \cbx_1__1_.Q_in[9] ;
 wire \cbx_1__1_.mux_bottom_ipin_0.INVTX1_4_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.INVTX1_5_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.INVTX1_3_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.INVTX1_4_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.INVTX1_5_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.INVTX1_3_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.INVTX1_5_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.INVTX1_3_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.INVTX1_4_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.INVTX1_5_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.INVTX1_3_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.INVTX1_4_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.INVTX1_5_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.INVTX1_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.INVTX1_3_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.INVTX1_4_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.INVTX1_5_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ;
 wire \cby_0__1_.Q_in[0] ;
 wire \cby_0__1_.Q_in[10] ;
 wire \cby_0__1_.Q_in[11] ;
 wire \cby_0__1_.Q_in[12] ;
 wire \cby_0__1_.Q_in[13] ;
 wire \cby_0__1_.Q_in[14] ;
 wire \cby_0__1_.Q_in[15] ;
 wire \cby_0__1_.Q_in[16] ;
 wire \cby_0__1_.Q_in[17] ;
 wire \cby_0__1_.Q_in[18] ;
 wire \cby_0__1_.Q_in[19] ;
 wire \cby_0__1_.Q_in[1] ;
 wire \cby_0__1_.Q_in[20] ;
 wire \cby_0__1_.Q_in[21] ;
 wire \cby_0__1_.Q_in[22] ;
 wire \cby_0__1_.Q_in[23] ;
 wire \cby_0__1_.Q_in[24] ;
 wire \cby_0__1_.Q_in[25] ;
 wire \cby_0__1_.Q_in[26] ;
 wire \cby_0__1_.Q_in[27] ;
 wire \cby_0__1_.Q_in[28] ;
 wire \cby_0__1_.Q_in[29] ;
 wire \cby_0__1_.Q_in[2] ;
 wire \cby_0__1_.Q_in[30] ;
 wire \cby_0__1_.Q_in[31] ;
 wire \cby_0__1_.Q_in[32] ;
 wire \cby_0__1_.Q_in[33] ;
 wire \cby_0__1_.Q_in[34] ;
 wire \cby_0__1_.Q_in[35] ;
 wire \cby_0__1_.Q_in[36] ;
 wire \cby_0__1_.Q_in[37] ;
 wire \cby_0__1_.Q_in[38] ;
 wire \cby_0__1_.Q_in[39] ;
 wire \cby_0__1_.Q_in[3] ;
 wire \cby_0__1_.Q_in[40] ;
 wire \cby_0__1_.Q_in[41] ;
 wire \cby_0__1_.Q_in[42] ;
 wire \cby_0__1_.Q_in[43] ;
 wire \cby_0__1_.Q_in[44] ;
 wire \cby_0__1_.Q_in[45] ;
 wire \cby_0__1_.Q_in[46] ;
 wire \cby_0__1_.Q_in[47] ;
 wire \cby_0__1_.Q_in[48] ;
 wire \cby_0__1_.Q_in[49] ;
 wire \cby_0__1_.Q_in[4] ;
 wire \cby_0__1_.Q_in[50] ;
 wire \cby_0__1_.Q_in[51] ;
 wire \cby_0__1_.Q_in[52] ;
 wire \cby_0__1_.Q_in[53] ;
 wire \cby_0__1_.Q_in[54] ;
 wire \cby_0__1_.Q_in[55] ;
 wire \cby_0__1_.Q_in[56] ;
 wire \cby_0__1_.Q_in[57] ;
 wire \cby_0__1_.Q_in[58] ;
 wire \cby_0__1_.Q_in[59] ;
 wire \cby_0__1_.Q_in[5] ;
 wire \cby_0__1_.Q_in[6] ;
 wire \cby_0__1_.Q_in[7] ;
 wire \cby_0__1_.Q_in[8] ;
 wire \cby_0__1_.Q_in[9] ;
 wire \cby_0__1_.mux_left_ipin_0.INVTX1_3_.out ;
 wire \cby_0__1_.mux_left_ipin_0.INVTX1_4_.out ;
 wire \cby_0__1_.mux_left_ipin_0.INVTX1_5_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ;
 wire \cby_0__1_.mux_left_ipin_1.INVTX1_2_.out ;
 wire \cby_0__1_.mux_left_ipin_1.INVTX1_4_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_0.INVTX1_2_.out ;
 wire \cby_0__1_.mux_right_ipin_0.INVTX1_3_.out ;
 wire \cby_0__1_.mux_right_ipin_0.INVTX1_4_.out ;
 wire \cby_0__1_.mux_right_ipin_0.INVTX1_5_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_1.INVTX1_2_.out ;
 wire \cby_0__1_.mux_right_ipin_1.INVTX1_3_.out ;
 wire \cby_0__1_.mux_right_ipin_1.INVTX1_5_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_2.INVTX1_2_.out ;
 wire \cby_0__1_.mux_right_ipin_2.INVTX1_3_.out ;
 wire \cby_0__1_.mux_right_ipin_2.INVTX1_5_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_3.INVTX1_2_.out ;
 wire \cby_0__1_.mux_right_ipin_3.INVTX1_3_.out ;
 wire \cby_0__1_.mux_right_ipin_3.INVTX1_4_.out ;
 wire \cby_0__1_.mux_right_ipin_3.INVTX1_5_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.Q_in[0] ;
 wire \cby_1__1_.Q_in[10] ;
 wire \cby_1__1_.Q_in[11] ;
 wire \cby_1__1_.Q_in[12] ;
 wire \cby_1__1_.Q_in[13] ;
 wire \cby_1__1_.Q_in[14] ;
 wire \cby_1__1_.Q_in[15] ;
 wire \cby_1__1_.Q_in[16] ;
 wire \cby_1__1_.Q_in[17] ;
 wire \cby_1__1_.Q_in[18] ;
 wire \cby_1__1_.Q_in[19] ;
 wire \cby_1__1_.Q_in[1] ;
 wire \cby_1__1_.Q_in[20] ;
 wire \cby_1__1_.Q_in[21] ;
 wire \cby_1__1_.Q_in[22] ;
 wire \cby_1__1_.Q_in[23] ;
 wire \cby_1__1_.Q_in[24] ;
 wire \cby_1__1_.Q_in[25] ;
 wire \cby_1__1_.Q_in[26] ;
 wire \cby_1__1_.Q_in[27] ;
 wire \cby_1__1_.Q_in[28] ;
 wire \cby_1__1_.Q_in[29] ;
 wire \cby_1__1_.Q_in[2] ;
 wire \cby_1__1_.Q_in[30] ;
 wire \cby_1__1_.Q_in[31] ;
 wire \cby_1__1_.Q_in[32] ;
 wire \cby_1__1_.Q_in[33] ;
 wire \cby_1__1_.Q_in[34] ;
 wire \cby_1__1_.Q_in[35] ;
 wire \cby_1__1_.Q_in[36] ;
 wire \cby_1__1_.Q_in[37] ;
 wire \cby_1__1_.Q_in[38] ;
 wire \cby_1__1_.Q_in[39] ;
 wire \cby_1__1_.Q_in[3] ;
 wire \cby_1__1_.Q_in[40] ;
 wire \cby_1__1_.Q_in[41] ;
 wire \cby_1__1_.Q_in[42] ;
 wire \cby_1__1_.Q_in[43] ;
 wire \cby_1__1_.Q_in[44] ;
 wire \cby_1__1_.Q_in[45] ;
 wire \cby_1__1_.Q_in[46] ;
 wire \cby_1__1_.Q_in[47] ;
 wire \cby_1__1_.Q_in[48] ;
 wire \cby_1__1_.Q_in[49] ;
 wire \cby_1__1_.Q_in[4] ;
 wire \cby_1__1_.Q_in[50] ;
 wire \cby_1__1_.Q_in[51] ;
 wire \cby_1__1_.Q_in[52] ;
 wire \cby_1__1_.Q_in[53] ;
 wire \cby_1__1_.Q_in[54] ;
 wire \cby_1__1_.Q_in[55] ;
 wire \cby_1__1_.Q_in[56] ;
 wire \cby_1__1_.Q_in[57] ;
 wire \cby_1__1_.Q_in[58] ;
 wire \cby_1__1_.Q_in[59] ;
 wire \cby_1__1_.Q_in[5] ;
 wire \cby_1__1_.Q_in[60] ;
 wire \cby_1__1_.Q_in[61] ;
 wire \cby_1__1_.Q_in[62] ;
 wire \cby_1__1_.Q_in[63] ;
 wire \cby_1__1_.Q_in[64] ;
 wire \cby_1__1_.Q_in[65] ;
 wire \cby_1__1_.Q_in[6] ;
 wire \cby_1__1_.Q_in[7] ;
 wire \cby_1__1_.Q_in[8] ;
 wire \cby_1__1_.Q_in[9] ;
 wire \cby_1__1_.mux_left_ipin_0.INVTX1_2_.out ;
 wire \cby_1__1_.mux_left_ipin_0.INVTX1_4_.out ;
 wire \cby_1__1_.mux_left_ipin_0.INVTX1_5_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_1.INVTX1_5_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_2.INVTX1_2_.out ;
 wire \cby_1__1_.mux_left_ipin_2.INVTX1_4_.out ;
 wire \cby_1__1_.mux_left_ipin_2.INVTX1_5_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_3.INVTX1_2_.out ;
 wire \cby_1__1_.mux_left_ipin_3.INVTX1_4_.out ;
 wire \cby_1__1_.mux_left_ipin_3.INVTX1_5_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_4.INVTX1_2_.out ;
 wire \cby_1__1_.mux_left_ipin_4.INVTX1_3_.out ;
 wire \cby_1__1_.mux_left_ipin_4.INVTX1_4_.out ;
 wire \cby_1__1_.mux_left_ipin_4.INVTX1_5_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_5.INVTX1_2_.out ;
 wire \cby_1__1_.mux_left_ipin_5.INVTX1_3_.out ;
 wire \cby_1__1_.mux_left_ipin_5.INVTX1_4_.out ;
 wire \cby_1__1_.mux_left_ipin_5.INVTX1_5_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ;
 wire \grid_clb_1__1_.Q_in[0] ;
 wire \grid_clb_1__1_.Q_in[100] ;
 wire \grid_clb_1__1_.Q_in[101] ;
 wire \grid_clb_1__1_.Q_in[102] ;
 wire \grid_clb_1__1_.Q_in[103] ;
 wire \grid_clb_1__1_.Q_in[104] ;
 wire \grid_clb_1__1_.Q_in[105] ;
 wire \grid_clb_1__1_.Q_in[106] ;
 wire \grid_clb_1__1_.Q_in[107] ;
 wire \grid_clb_1__1_.Q_in[108] ;
 wire \grid_clb_1__1_.Q_in[109] ;
 wire \grid_clb_1__1_.Q_in[10] ;
 wire \grid_clb_1__1_.Q_in[110] ;
 wire \grid_clb_1__1_.Q_in[111] ;
 wire \grid_clb_1__1_.Q_in[112] ;
 wire \grid_clb_1__1_.Q_in[113] ;
 wire \grid_clb_1__1_.Q_in[114] ;
 wire \grid_clb_1__1_.Q_in[115] ;
 wire \grid_clb_1__1_.Q_in[116] ;
 wire \grid_clb_1__1_.Q_in[117] ;
 wire \grid_clb_1__1_.Q_in[118] ;
 wire \grid_clb_1__1_.Q_in[119] ;
 wire \grid_clb_1__1_.Q_in[11] ;
 wire \grid_clb_1__1_.Q_in[120] ;
 wire \grid_clb_1__1_.Q_in[121] ;
 wire \grid_clb_1__1_.Q_in[122] ;
 wire \grid_clb_1__1_.Q_in[123] ;
 wire \grid_clb_1__1_.Q_in[124] ;
 wire \grid_clb_1__1_.Q_in[125] ;
 wire \grid_clb_1__1_.Q_in[126] ;
 wire \grid_clb_1__1_.Q_in[127] ;
 wire \grid_clb_1__1_.Q_in[128] ;
 wire \grid_clb_1__1_.Q_in[129] ;
 wire \grid_clb_1__1_.Q_in[12] ;
 wire \grid_clb_1__1_.Q_in[130] ;
 wire \grid_clb_1__1_.Q_in[131] ;
 wire \grid_clb_1__1_.Q_in[132] ;
 wire \grid_clb_1__1_.Q_in[133] ;
 wire \grid_clb_1__1_.Q_in[134] ;
 wire \grid_clb_1__1_.Q_in[135] ;
 wire \grid_clb_1__1_.Q_in[136] ;
 wire \grid_clb_1__1_.Q_in[137] ;
 wire \grid_clb_1__1_.Q_in[138] ;
 wire \grid_clb_1__1_.Q_in[139] ;
 wire \grid_clb_1__1_.Q_in[13] ;
 wire \grid_clb_1__1_.Q_in[140] ;
 wire \grid_clb_1__1_.Q_in[141] ;
 wire \grid_clb_1__1_.Q_in[142] ;
 wire \grid_clb_1__1_.Q_in[143] ;
 wire \grid_clb_1__1_.Q_in[144] ;
 wire \grid_clb_1__1_.Q_in[145] ;
 wire \grid_clb_1__1_.Q_in[146] ;
 wire \grid_clb_1__1_.Q_in[147] ;
 wire \grid_clb_1__1_.Q_in[148] ;
 wire \grid_clb_1__1_.Q_in[149] ;
 wire \grid_clb_1__1_.Q_in[14] ;
 wire \grid_clb_1__1_.Q_in[150] ;
 wire \grid_clb_1__1_.Q_in[151] ;
 wire \grid_clb_1__1_.Q_in[152] ;
 wire \grid_clb_1__1_.Q_in[153] ;
 wire \grid_clb_1__1_.Q_in[154] ;
 wire \grid_clb_1__1_.Q_in[155] ;
 wire \grid_clb_1__1_.Q_in[156] ;
 wire \grid_clb_1__1_.Q_in[157] ;
 wire \grid_clb_1__1_.Q_in[158] ;
 wire \grid_clb_1__1_.Q_in[159] ;
 wire \grid_clb_1__1_.Q_in[15] ;
 wire \grid_clb_1__1_.Q_in[160] ;
 wire \grid_clb_1__1_.Q_in[161] ;
 wire \grid_clb_1__1_.Q_in[162] ;
 wire \grid_clb_1__1_.Q_in[163] ;
 wire \grid_clb_1__1_.Q_in[164] ;
 wire \grid_clb_1__1_.Q_in[165] ;
 wire \grid_clb_1__1_.Q_in[166] ;
 wire \grid_clb_1__1_.Q_in[167] ;
 wire \grid_clb_1__1_.Q_in[168] ;
 wire \grid_clb_1__1_.Q_in[169] ;
 wire \grid_clb_1__1_.Q_in[16] ;
 wire \grid_clb_1__1_.Q_in[170] ;
 wire \grid_clb_1__1_.Q_in[171] ;
 wire \grid_clb_1__1_.Q_in[172] ;
 wire \grid_clb_1__1_.Q_in[173] ;
 wire \grid_clb_1__1_.Q_in[174] ;
 wire \grid_clb_1__1_.Q_in[175] ;
 wire \grid_clb_1__1_.Q_in[176] ;
 wire \grid_clb_1__1_.Q_in[177] ;
 wire \grid_clb_1__1_.Q_in[178] ;
 wire \grid_clb_1__1_.Q_in[179] ;
 wire \grid_clb_1__1_.Q_in[17] ;
 wire \grid_clb_1__1_.Q_in[180] ;
 wire \grid_clb_1__1_.Q_in[181] ;
 wire \grid_clb_1__1_.Q_in[182] ;
 wire \grid_clb_1__1_.Q_in[183] ;
 wire \grid_clb_1__1_.Q_in[184] ;
 wire \grid_clb_1__1_.Q_in[185] ;
 wire \grid_clb_1__1_.Q_in[186] ;
 wire \grid_clb_1__1_.Q_in[187] ;
 wire \grid_clb_1__1_.Q_in[188] ;
 wire \grid_clb_1__1_.Q_in[189] ;
 wire \grid_clb_1__1_.Q_in[18] ;
 wire \grid_clb_1__1_.Q_in[190] ;
 wire \grid_clb_1__1_.Q_in[191] ;
 wire \grid_clb_1__1_.Q_in[192] ;
 wire \grid_clb_1__1_.Q_in[193] ;
 wire \grid_clb_1__1_.Q_in[194] ;
 wire \grid_clb_1__1_.Q_in[195] ;
 wire \grid_clb_1__1_.Q_in[196] ;
 wire \grid_clb_1__1_.Q_in[197] ;
 wire \grid_clb_1__1_.Q_in[198] ;
 wire \grid_clb_1__1_.Q_in[199] ;
 wire \grid_clb_1__1_.Q_in[19] ;
 wire \grid_clb_1__1_.Q_in[1] ;
 wire \grid_clb_1__1_.Q_in[200] ;
 wire \grid_clb_1__1_.Q_in[201] ;
 wire \grid_clb_1__1_.Q_in[202] ;
 wire \grid_clb_1__1_.Q_in[203] ;
 wire \grid_clb_1__1_.Q_in[20] ;
 wire \grid_clb_1__1_.Q_in[21] ;
 wire \grid_clb_1__1_.Q_in[22] ;
 wire \grid_clb_1__1_.Q_in[23] ;
 wire \grid_clb_1__1_.Q_in[24] ;
 wire \grid_clb_1__1_.Q_in[25] ;
 wire \grid_clb_1__1_.Q_in[26] ;
 wire \grid_clb_1__1_.Q_in[27] ;
 wire \grid_clb_1__1_.Q_in[28] ;
 wire \grid_clb_1__1_.Q_in[29] ;
 wire \grid_clb_1__1_.Q_in[2] ;
 wire \grid_clb_1__1_.Q_in[30] ;
 wire \grid_clb_1__1_.Q_in[31] ;
 wire \grid_clb_1__1_.Q_in[32] ;
 wire \grid_clb_1__1_.Q_in[33] ;
 wire \grid_clb_1__1_.Q_in[34] ;
 wire \grid_clb_1__1_.Q_in[35] ;
 wire \grid_clb_1__1_.Q_in[36] ;
 wire \grid_clb_1__1_.Q_in[37] ;
 wire \grid_clb_1__1_.Q_in[38] ;
 wire \grid_clb_1__1_.Q_in[39] ;
 wire \grid_clb_1__1_.Q_in[3] ;
 wire \grid_clb_1__1_.Q_in[40] ;
 wire \grid_clb_1__1_.Q_in[41] ;
 wire \grid_clb_1__1_.Q_in[42] ;
 wire \grid_clb_1__1_.Q_in[43] ;
 wire \grid_clb_1__1_.Q_in[44] ;
 wire \grid_clb_1__1_.Q_in[45] ;
 wire \grid_clb_1__1_.Q_in[46] ;
 wire \grid_clb_1__1_.Q_in[47] ;
 wire \grid_clb_1__1_.Q_in[48] ;
 wire \grid_clb_1__1_.Q_in[49] ;
 wire \grid_clb_1__1_.Q_in[4] ;
 wire \grid_clb_1__1_.Q_in[50] ;
 wire \grid_clb_1__1_.Q_in[51] ;
 wire \grid_clb_1__1_.Q_in[52] ;
 wire \grid_clb_1__1_.Q_in[53] ;
 wire \grid_clb_1__1_.Q_in[54] ;
 wire \grid_clb_1__1_.Q_in[55] ;
 wire \grid_clb_1__1_.Q_in[56] ;
 wire \grid_clb_1__1_.Q_in[57] ;
 wire \grid_clb_1__1_.Q_in[58] ;
 wire \grid_clb_1__1_.Q_in[59] ;
 wire \grid_clb_1__1_.Q_in[5] ;
 wire \grid_clb_1__1_.Q_in[60] ;
 wire \grid_clb_1__1_.Q_in[61] ;
 wire \grid_clb_1__1_.Q_in[62] ;
 wire \grid_clb_1__1_.Q_in[63] ;
 wire \grid_clb_1__1_.Q_in[64] ;
 wire \grid_clb_1__1_.Q_in[65] ;
 wire \grid_clb_1__1_.Q_in[66] ;
 wire \grid_clb_1__1_.Q_in[67] ;
 wire \grid_clb_1__1_.Q_in[68] ;
 wire \grid_clb_1__1_.Q_in[69] ;
 wire \grid_clb_1__1_.Q_in[6] ;
 wire \grid_clb_1__1_.Q_in[70] ;
 wire \grid_clb_1__1_.Q_in[71] ;
 wire \grid_clb_1__1_.Q_in[72] ;
 wire \grid_clb_1__1_.Q_in[73] ;
 wire \grid_clb_1__1_.Q_in[74] ;
 wire \grid_clb_1__1_.Q_in[75] ;
 wire \grid_clb_1__1_.Q_in[76] ;
 wire \grid_clb_1__1_.Q_in[77] ;
 wire \grid_clb_1__1_.Q_in[78] ;
 wire \grid_clb_1__1_.Q_in[79] ;
 wire \grid_clb_1__1_.Q_in[7] ;
 wire \grid_clb_1__1_.Q_in[80] ;
 wire \grid_clb_1__1_.Q_in[81] ;
 wire \grid_clb_1__1_.Q_in[82] ;
 wire \grid_clb_1__1_.Q_in[83] ;
 wire \grid_clb_1__1_.Q_in[84] ;
 wire \grid_clb_1__1_.Q_in[85] ;
 wire \grid_clb_1__1_.Q_in[86] ;
 wire \grid_clb_1__1_.Q_in[87] ;
 wire \grid_clb_1__1_.Q_in[88] ;
 wire \grid_clb_1__1_.Q_in[89] ;
 wire \grid_clb_1__1_.Q_in[8] ;
 wire \grid_clb_1__1_.Q_in[90] ;
 wire \grid_clb_1__1_.Q_in[91] ;
 wire \grid_clb_1__1_.Q_in[92] ;
 wire \grid_clb_1__1_.Q_in[93] ;
 wire \grid_clb_1__1_.Q_in[94] ;
 wire \grid_clb_1__1_.Q_in[95] ;
 wire \grid_clb_1__1_.Q_in[96] ;
 wire \grid_clb_1__1_.Q_in[97] ;
 wire \grid_clb_1__1_.Q_in[98] ;
 wire \grid_clb_1__1_.Q_in[99] ;
 wire \grid_clb_1__1_.Q_in[9] ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_ff_0.DFFSRQ_0_.D ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_ff_0.DFFSRQ_0_.D ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_ff_0.DFFSRQ_0_.D ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_ff_0.DFFSRQ_0_.D ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.INVTX1_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.out ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[0] ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[1] ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[2] ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[3] ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[4] ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[5] ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[6] ;
 wire \grid_io_bottom_1__0_.GPIO_DIR[7] ;
 wire \grid_io_left_0__1_.GPIO_DIR[0] ;
 wire \grid_io_left_0__1_.GPIO_DIR[1] ;
 wire \grid_io_left_0__1_.GPIO_DIR[2] ;
 wire \grid_io_left_0__1_.GPIO_DIR[3] ;
 wire \grid_io_left_0__1_.GPIO_DIR[4] ;
 wire \grid_io_left_0__1_.GPIO_DIR[5] ;
 wire \grid_io_left_0__1_.GPIO_DIR[6] ;
 wire \grid_io_left_0__1_.GPIO_DIR[7] ;
 wire \grid_io_right_2__1_.GPIO_DIR[0] ;
 wire \grid_io_right_2__1_.GPIO_DIR[1] ;
 wire \grid_io_right_2__1_.GPIO_DIR[2] ;
 wire \grid_io_right_2__1_.GPIO_DIR[3] ;
 wire \grid_io_right_2__1_.GPIO_DIR[4] ;
 wire \grid_io_right_2__1_.GPIO_DIR[5] ;
 wire \grid_io_right_2__1_.GPIO_DIR[6] ;
 wire \grid_io_right_2__1_.GPIO_DIR[7] ;
 wire \grid_io_top_1__2_.GPIO_DIR[0] ;
 wire \grid_io_top_1__2_.GPIO_DIR[1] ;
 wire \grid_io_top_1__2_.GPIO_DIR[2] ;
 wire \grid_io_top_1__2_.GPIO_DIR[3] ;
 wire \grid_io_top_1__2_.GPIO_DIR[4] ;
 wire \grid_io_top_1__2_.GPIO_DIR[5] ;
 wire \grid_io_top_1__2_.GPIO_DIR[6] ;
 wire \grid_io_top_1__2_.GPIO_DIR[7] ;
 wire \sb_0__0_.Q_in[0] ;
 wire \sb_0__0_.Q_in[10] ;
 wire \sb_0__0_.Q_in[11] ;
 wire \sb_0__0_.Q_in[12] ;
 wire \sb_0__0_.Q_in[13] ;
 wire \sb_0__0_.Q_in[14] ;
 wire \sb_0__0_.Q_in[15] ;
 wire \sb_0__0_.Q_in[16] ;
 wire \sb_0__0_.Q_in[17] ;
 wire \sb_0__0_.Q_in[18] ;
 wire \sb_0__0_.Q_in[19] ;
 wire \sb_0__0_.Q_in[1] ;
 wire \sb_0__0_.Q_in[20] ;
 wire \sb_0__0_.Q_in[21] ;
 wire \sb_0__0_.Q_in[22] ;
 wire \sb_0__0_.Q_in[23] ;
 wire \sb_0__0_.Q_in[24] ;
 wire \sb_0__0_.Q_in[25] ;
 wire \sb_0__0_.Q_in[26] ;
 wire \sb_0__0_.Q_in[27] ;
 wire \sb_0__0_.Q_in[28] ;
 wire \sb_0__0_.Q_in[29] ;
 wire \sb_0__0_.Q_in[2] ;
 wire \sb_0__0_.Q_in[30] ;
 wire \sb_0__0_.Q_in[31] ;
 wire \sb_0__0_.Q_in[32] ;
 wire \sb_0__0_.Q_in[33] ;
 wire \sb_0__0_.Q_in[34] ;
 wire \sb_0__0_.Q_in[35] ;
 wire \sb_0__0_.Q_in[36] ;
 wire \sb_0__0_.Q_in[37] ;
 wire \sb_0__0_.Q_in[38] ;
 wire \sb_0__0_.Q_in[39] ;
 wire \sb_0__0_.Q_in[3] ;
 wire \sb_0__0_.Q_in[40] ;
 wire \sb_0__0_.Q_in[41] ;
 wire \sb_0__0_.Q_in[42] ;
 wire \sb_0__0_.Q_in[43] ;
 wire \sb_0__0_.Q_in[44] ;
 wire \sb_0__0_.Q_in[45] ;
 wire \sb_0__0_.Q_in[46] ;
 wire \sb_0__0_.Q_in[47] ;
 wire \sb_0__0_.Q_in[48] ;
 wire \sb_0__0_.Q_in[49] ;
 wire \sb_0__0_.Q_in[4] ;
 wire \sb_0__0_.Q_in[50] ;
 wire \sb_0__0_.Q_in[51] ;
 wire \sb_0__0_.Q_in[52] ;
 wire \sb_0__0_.Q_in[53] ;
 wire \sb_0__0_.Q_in[54] ;
 wire \sb_0__0_.Q_in[55] ;
 wire \sb_0__0_.Q_in[56] ;
 wire \sb_0__0_.Q_in[57] ;
 wire \sb_0__0_.Q_in[58] ;
 wire \sb_0__0_.Q_in[59] ;
 wire \sb_0__0_.Q_in[5] ;
 wire \sb_0__0_.Q_in[60] ;
 wire \sb_0__0_.Q_in[61] ;
 wire \sb_0__0_.Q_in[62] ;
 wire \sb_0__0_.Q_in[63] ;
 wire \sb_0__0_.Q_in[64] ;
 wire \sb_0__0_.Q_in[65] ;
 wire \sb_0__0_.Q_in[66] ;
 wire \sb_0__0_.Q_in[67] ;
 wire \sb_0__0_.Q_in[68] ;
 wire \sb_0__0_.Q_in[69] ;
 wire \sb_0__0_.Q_in[6] ;
 wire \sb_0__0_.Q_in[70] ;
 wire \sb_0__0_.Q_in[71] ;
 wire \sb_0__0_.Q_in[72] ;
 wire \sb_0__0_.Q_in[73] ;
 wire \sb_0__0_.Q_in[74] ;
 wire \sb_0__0_.Q_in[75] ;
 wire \sb_0__0_.Q_in[7] ;
 wire \sb_0__0_.Q_in[8] ;
 wire \sb_0__0_.Q_in[9] ;
 wire \sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_0.mux_l1_in_0_.out ;
 wire \sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_0.mux_l2_in_0_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l1_in_0_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_12.mux_l2_in_0_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l1_in_0_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_14.mux_l2_in_0_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l1_in_0_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_right_track_2.mux_l2_in_0_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l1_in_0_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_top_track_0.mux_l2_in_0_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l1_in_0_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__0_.mux_top_track_12.mux_l2_in_0_.out ;
 wire \sb_0__1_.Q_in[14] ;
 wire \sb_0__1_.Q_in[15] ;
 wire \sb_0__1_.Q_in[16] ;
 wire \sb_0__1_.Q_in[17] ;
 wire \sb_0__1_.Q_in[18] ;
 wire \sb_0__1_.Q_in[19] ;
 wire \sb_0__1_.Q_in[20] ;
 wire \sb_0__1_.Q_in[21] ;
 wire \sb_0__1_.Q_in[22] ;
 wire \sb_0__1_.Q_in[23] ;
 wire \sb_0__1_.Q_in[24] ;
 wire \sb_0__1_.Q_in[25] ;
 wire \sb_0__1_.Q_in[26] ;
 wire \sb_0__1_.Q_in[27] ;
 wire \sb_0__1_.Q_in[28] ;
 wire \sb_0__1_.Q_in[29] ;
 wire \sb_0__1_.Q_in[30] ;
 wire \sb_0__1_.Q_in[31] ;
 wire \sb_0__1_.Q_in[32] ;
 wire \sb_0__1_.Q_in[33] ;
 wire \sb_0__1_.Q_in[34] ;
 wire \sb_0__1_.Q_in[35] ;
 wire \sb_0__1_.Q_in[36] ;
 wire \sb_0__1_.Q_in[37] ;
 wire \sb_0__1_.Q_in[38] ;
 wire \sb_0__1_.Q_in[39] ;
 wire \sb_0__1_.Q_in[40] ;
 wire \sb_0__1_.Q_in[41] ;
 wire \sb_0__1_.Q_in[42] ;
 wire \sb_0__1_.Q_in[43] ;
 wire \sb_0__1_.Q_in[44] ;
 wire \sb_0__1_.Q_in[45] ;
 wire \sb_0__1_.Q_in[46] ;
 wire \sb_0__1_.Q_in[47] ;
 wire \sb_0__1_.Q_in[48] ;
 wire \sb_0__1_.Q_in[49] ;
 wire \sb_0__1_.Q_in[50] ;
 wire \sb_0__1_.Q_in[51] ;
 wire \sb_0__1_.Q_in[52] ;
 wire \sb_0__1_.Q_in[53] ;
 wire \sb_0__1_.Q_in[54] ;
 wire \sb_0__1_.Q_in[55] ;
 wire \sb_0__1_.Q_in[56] ;
 wire \sb_0__1_.Q_in[57] ;
 wire \sb_0__1_.Q_in[58] ;
 wire \sb_0__1_.Q_in[59] ;
 wire \sb_0__1_.Q_in[60] ;
 wire \sb_0__1_.Q_in[61] ;
 wire \sb_0__1_.Q_in[62] ;
 wire \sb_0__1_.Q_in[63] ;
 wire \sb_0__1_.Q_in[64] ;
 wire \sb_0__1_.Q_in[65] ;
 wire \sb_0__1_.Q_in[66] ;
 wire \sb_0__1_.Q_in[67] ;
 wire \sb_0__1_.Q_in[68] ;
 wire \sb_0__1_.Q_in[69] ;
 wire \sb_0__1_.Q_in[70] ;
 wire \sb_0__1_.Q_in[71] ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.out ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l1_in_0_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_right_track_0.mux_l2_in_0_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l1_in_0_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_0__1_.mux_right_track_12.mux_l2_in_0_.out ;
 wire \sb_1__0_.Q_in[0] ;
 wire \sb_1__0_.Q_in[10] ;
 wire \sb_1__0_.Q_in[11] ;
 wire \sb_1__0_.Q_in[12] ;
 wire \sb_1__0_.Q_in[13] ;
 wire \sb_1__0_.Q_in[14] ;
 wire \sb_1__0_.Q_in[15] ;
 wire \sb_1__0_.Q_in[16] ;
 wire \sb_1__0_.Q_in[17] ;
 wire \sb_1__0_.Q_in[18] ;
 wire \sb_1__0_.Q_in[19] ;
 wire \sb_1__0_.Q_in[1] ;
 wire \sb_1__0_.Q_in[20] ;
 wire \sb_1__0_.Q_in[21] ;
 wire \sb_1__0_.Q_in[22] ;
 wire \sb_1__0_.Q_in[23] ;
 wire \sb_1__0_.Q_in[24] ;
 wire \sb_1__0_.Q_in[25] ;
 wire \sb_1__0_.Q_in[26] ;
 wire \sb_1__0_.Q_in[27] ;
 wire \sb_1__0_.Q_in[28] ;
 wire \sb_1__0_.Q_in[29] ;
 wire \sb_1__0_.Q_in[2] ;
 wire \sb_1__0_.Q_in[30] ;
 wire \sb_1__0_.Q_in[31] ;
 wire \sb_1__0_.Q_in[32] ;
 wire \sb_1__0_.Q_in[33] ;
 wire \sb_1__0_.Q_in[34] ;
 wire \sb_1__0_.Q_in[35] ;
 wire \sb_1__0_.Q_in[36] ;
 wire \sb_1__0_.Q_in[37] ;
 wire \sb_1__0_.Q_in[38] ;
 wire \sb_1__0_.Q_in[39] ;
 wire \sb_1__0_.Q_in[3] ;
 wire \sb_1__0_.Q_in[40] ;
 wire \sb_1__0_.Q_in[41] ;
 wire \sb_1__0_.Q_in[42] ;
 wire \sb_1__0_.Q_in[43] ;
 wire \sb_1__0_.Q_in[44] ;
 wire \sb_1__0_.Q_in[45] ;
 wire \sb_1__0_.Q_in[46] ;
 wire \sb_1__0_.Q_in[47] ;
 wire \sb_1__0_.Q_in[48] ;
 wire \sb_1__0_.Q_in[49] ;
 wire \sb_1__0_.Q_in[4] ;
 wire \sb_1__0_.Q_in[50] ;
 wire \sb_1__0_.Q_in[51] ;
 wire \sb_1__0_.Q_in[52] ;
 wire \sb_1__0_.Q_in[53] ;
 wire \sb_1__0_.Q_in[54] ;
 wire \sb_1__0_.Q_in[55] ;
 wire \sb_1__0_.Q_in[56] ;
 wire \sb_1__0_.Q_in[57] ;
 wire \sb_1__0_.Q_in[58] ;
 wire \sb_1__0_.Q_in[59] ;
 wire \sb_1__0_.Q_in[5] ;
 wire \sb_1__0_.Q_in[60] ;
 wire \sb_1__0_.Q_in[61] ;
 wire \sb_1__0_.Q_in[62] ;
 wire \sb_1__0_.Q_in[63] ;
 wire \sb_1__0_.Q_in[64] ;
 wire \sb_1__0_.Q_in[65] ;
 wire \sb_1__0_.Q_in[66] ;
 wire \sb_1__0_.Q_in[67] ;
 wire \sb_1__0_.Q_in[68] ;
 wire \sb_1__0_.Q_in[69] ;
 wire \sb_1__0_.Q_in[6] ;
 wire \sb_1__0_.Q_in[70] ;
 wire \sb_1__0_.Q_in[71] ;
 wire \sb_1__0_.Q_in[72] ;
 wire \sb_1__0_.Q_in[73] ;
 wire \sb_1__0_.Q_in[74] ;
 wire \sb_1__0_.Q_in[75] ;
 wire \sb_1__0_.Q_in[76] ;
 wire \sb_1__0_.Q_in[77] ;
 wire \sb_1__0_.Q_in[78] ;
 wire \sb_1__0_.Q_in[79] ;
 wire \sb_1__0_.Q_in[7] ;
 wire \sb_1__0_.Q_in[8] ;
 wire \sb_1__0_.Q_in[9] ;
 wire \sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_1.mux_l1_in_0_.out ;
 wire \sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_1.mux_l2_in_0_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l1_in_0_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_13.mux_l2_in_0_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l1_in_0_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_15.mux_l2_in_0_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l1_in_0_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_left_track_3.mux_l2_in_0_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l1_in_0_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l1_in_0_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_top_track_14.mux_l2_in_0_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l1_in_0_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__0_.mux_top_track_2.mux_l2_in_0_.out ;
 wire \sb_1__1_.Q_in[0] ;
 wire \sb_1__1_.Q_in[10] ;
 wire \sb_1__1_.Q_in[11] ;
 wire \sb_1__1_.Q_in[12] ;
 wire \sb_1__1_.Q_in[13] ;
 wire \sb_1__1_.Q_in[14] ;
 wire \sb_1__1_.Q_in[15] ;
 wire \sb_1__1_.Q_in[16] ;
 wire \sb_1__1_.Q_in[17] ;
 wire \sb_1__1_.Q_in[18] ;
 wire \sb_1__1_.Q_in[19] ;
 wire \sb_1__1_.Q_in[1] ;
 wire \sb_1__1_.Q_in[20] ;
 wire \sb_1__1_.Q_in[21] ;
 wire \sb_1__1_.Q_in[22] ;
 wire \sb_1__1_.Q_in[23] ;
 wire \sb_1__1_.Q_in[24] ;
 wire \sb_1__1_.Q_in[25] ;
 wire \sb_1__1_.Q_in[26] ;
 wire \sb_1__1_.Q_in[27] ;
 wire \sb_1__1_.Q_in[28] ;
 wire \sb_1__1_.Q_in[29] ;
 wire \sb_1__1_.Q_in[2] ;
 wire \sb_1__1_.Q_in[30] ;
 wire \sb_1__1_.Q_in[31] ;
 wire \sb_1__1_.Q_in[32] ;
 wire \sb_1__1_.Q_in[33] ;
 wire \sb_1__1_.Q_in[34] ;
 wire \sb_1__1_.Q_in[35] ;
 wire \sb_1__1_.Q_in[36] ;
 wire \sb_1__1_.Q_in[37] ;
 wire \sb_1__1_.Q_in[38] ;
 wire \sb_1__1_.Q_in[39] ;
 wire \sb_1__1_.Q_in[3] ;
 wire \sb_1__1_.Q_in[40] ;
 wire \sb_1__1_.Q_in[41] ;
 wire \sb_1__1_.Q_in[42] ;
 wire \sb_1__1_.Q_in[43] ;
 wire \sb_1__1_.Q_in[44] ;
 wire \sb_1__1_.Q_in[45] ;
 wire \sb_1__1_.Q_in[46] ;
 wire \sb_1__1_.Q_in[47] ;
 wire \sb_1__1_.Q_in[48] ;
 wire \sb_1__1_.Q_in[49] ;
 wire \sb_1__1_.Q_in[4] ;
 wire \sb_1__1_.Q_in[50] ;
 wire \sb_1__1_.Q_in[51] ;
 wire \sb_1__1_.Q_in[52] ;
 wire \sb_1__1_.Q_in[53] ;
 wire \sb_1__1_.Q_in[54] ;
 wire \sb_1__1_.Q_in[55] ;
 wire \sb_1__1_.Q_in[56] ;
 wire \sb_1__1_.Q_in[57] ;
 wire \sb_1__1_.Q_in[58] ;
 wire \sb_1__1_.Q_in[59] ;
 wire \sb_1__1_.Q_in[5] ;
 wire \sb_1__1_.Q_in[60] ;
 wire \sb_1__1_.Q_in[61] ;
 wire \sb_1__1_.Q_in[62] ;
 wire \sb_1__1_.Q_in[63] ;
 wire \sb_1__1_.Q_in[64] ;
 wire \sb_1__1_.Q_in[65] ;
 wire \sb_1__1_.Q_in[66] ;
 wire \sb_1__1_.Q_in[67] ;
 wire \sb_1__1_.Q_in[6] ;
 wire \sb_1__1_.Q_in[7] ;
 wire \sb_1__1_.Q_in[8] ;
 wire \sb_1__1_.Q_in[9] ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.out ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l1_in_0_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_left_track_1.mux_l2_in_0_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l1_in_0_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.out ;
 wire \sb_1__1_.mux_left_track_13.mux_l2_in_0_.out ;

 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_590 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_96 ();
 sky130_fd_sc_hd__or3_1 _0726_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0727_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0728_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0729_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0730_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0731_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0732_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0733_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0734_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0735_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0736_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0737_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0738_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0739_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0740_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0741_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0742_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0743_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0744_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0745_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0746_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0747_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0748_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0749_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0750_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0751_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0752_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0753_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0754_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0755_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0756_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0757_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0758_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0759_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0760_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0761_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0762_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0763_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0764_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0765_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0766_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0767_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0768_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0769_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0770_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0771_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0772_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0773_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0774_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0775_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0776_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0777_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0778_ (.A(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0779_ (.A(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0780_ (.A(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0781_ (.A(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0782_ (.A(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0783_ (.A(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0784_ (.A(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0785_ (.A(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0786_ (.A(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0787_ (.A(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0788_ (.A(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0789_ (.A(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0790_ (.A(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_1 _0791_ (.A(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.out ),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_1 _0792_ (.A(_0520_),
    .Y(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0793_ (.A(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_1 _0794_ (.A(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.out ),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_1 _0795_ (.A(_0521_),
    .Y(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0796_ (.A(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0797_ (.A(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0798_ (.A(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0799_ (.A(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0800_ (.A(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0801_ (.A(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0802_ (.A(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0803_ (.A(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0804_ (.A(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0805_ (.A(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0806_ (.A(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0807_ (.A(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0808_ (.A(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_2 _0809_ (.A(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_1 _0810_ (.A(_0522_),
    .Y(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0811_ (.A(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0812_ (.A(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0813_ (.A(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_1 _0814_ (.A(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.out ),
    .Y(_0523_));
 sky130_fd_sc_hd__inv_1 _0815_ (.A(_0523_),
    .Y(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0816_ (.A(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_4 _0817_ (.A(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0818_ (.A(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_1 _0819_ (.A(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.out ),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_1 _0820_ (.A(_0524_),
    .Y(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0821_ (.A(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_1 _0822_ (.A(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_1 _0823_ (.A(_0525_),
    .Y(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0824_ (.A(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0825_ (.A(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0826_ (.A(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0827_ (.A(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ),
    .X(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0828_ (.A(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0829_ (.A(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0830_ (.A(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0831_ (.A(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0832_ (.A(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0833_ (.A(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0834_ (.A(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0835_ (.A(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0836_ (.A(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0837_ (.A(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0838_ (.A(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0839_ (.A(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0840_ (.A(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0841_ (.A(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0842_ (.A(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0843_ (.A(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0844_ (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0845_ (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0846_ (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0847_ (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0848_ (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0849_ (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0850_ (.A(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0851_ (.A(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0852_ (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0853_ (.A(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0854_ (.A(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0855_ (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0856_ (.A(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0857_ (.A(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0858_ (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0859_ (.A(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0860_ (.A(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0861_ (.A(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0862_ (.A(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0863_ (.A(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0864_ (.A(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0865_ (.A(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0866_ (.A(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0867_ (.A(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0868_ (.A(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0869_ (.A(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0870_ (.A(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0871_ (.A(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0872_ (.A(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0873_ (.A(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0874_ (.A(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0875_ (.A(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0876_ (.A(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0877_ (.A(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0878_ (.A(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0879_ (.A(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0880_ (.A(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0881_ (.A(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0882_ (.A(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0883_ (.A(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0884_ (.A(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0885_ (.A(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0886_ (.A(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0887_ (.A(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0888_ (.A(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0889_ (.A(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0890_ (.A(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0891_ (.A(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0892_ (.A(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0893_ (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0894_ (.A(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0895_ (.A(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0896_ (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0897_ (.A(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0898_ (.A(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0899_ (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0900_ (.A(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0901_ (.A(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0902_ (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0903_ (.A(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0904_ (.A(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0905_ (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0906_ (.A(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0907_ (.A(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0908_ (.A(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0909_ (.A(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0910_ (.A(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0911_ (.A(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0912_ (.A(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0913_ (.A(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0914_ (.A(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0915_ (.A(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0916_ (.A(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0917_ (.A(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0918_ (.A(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0919_ (.A(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0920_ (.A(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0921_ (.A(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out ),
    .X(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or3_1 _0922_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_1 _0923_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_1 _0924_ (.A(_0526_),
    .Y(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0925_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor3_1 _0926_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ),
    .Y(_0527_));
 sky130_fd_sc_hd__inv_1 _0927_ (.A(_0527_),
    .Y(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0928_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0929_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0930_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0931_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0932_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0933_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0934_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0935_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__or3_1 _0936_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.out ));
 sky130_fd_sc_hd__or4_1 _0937_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.out ));
 sky130_fd_sc_hd__or4_1 _0938_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.out ));
 sky130_fd_sc_hd__or4_1 _0939_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.out ),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.out ));
 sky130_fd_sc_hd__nor4_1 _0940_ (.A(\cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[7] ),
    .Y(gfpga_pad_GPIO_PAD[7]));
 sky130_fd_sc_hd__nor4_1 _0941_ (.A(\cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[6] ),
    .Y(gfpga_pad_GPIO_PAD[6]));
 sky130_fd_sc_hd__nor4_1 _0942_ (.A(\cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[5] ),
    .Y(gfpga_pad_GPIO_PAD[5]));
 sky130_fd_sc_hd__nor4_1 _0943_ (.A(\cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[4] ),
    .Y(gfpga_pad_GPIO_PAD[4]));
 sky130_fd_sc_hd__nor4_1 _0944_ (.A(\cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[3] ),
    .Y(gfpga_pad_GPIO_PAD[3]));
 sky130_fd_sc_hd__nor4_1 _0945_ (.A(\cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[2] ),
    .Y(gfpga_pad_GPIO_PAD[2]));
 sky130_fd_sc_hd__nor4_1 _0946_ (.A(\cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[1] ),
    .Y(gfpga_pad_GPIO_PAD[1]));
 sky130_fd_sc_hd__nor4_1 _0947_ (.A(\cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_top_1__2_.GPIO_DIR[0] ),
    .Y(gfpga_pad_GPIO_PAD[0]));
 sky130_fd_sc_hd__nor4_1 _0948_ (.A(\cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[7] ),
    .Y(gfpga_pad_GPIO_PAD[15]));
 sky130_fd_sc_hd__nor4_1 _0949_ (.A(\cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[6] ),
    .Y(gfpga_pad_GPIO_PAD[14]));
 sky130_fd_sc_hd__nor4_1 _0950_ (.A(\cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[5] ),
    .Y(gfpga_pad_GPIO_PAD[13]));
 sky130_fd_sc_hd__nor4_1 _0951_ (.A(\cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[4] ),
    .Y(gfpga_pad_GPIO_PAD[12]));
 sky130_fd_sc_hd__nor4_1 _0952_ (.A(\cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[3] ),
    .Y(gfpga_pad_GPIO_PAD[11]));
 sky130_fd_sc_hd__nor4_1 _0953_ (.A(\cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[2] ),
    .Y(gfpga_pad_GPIO_PAD[10]));
 sky130_fd_sc_hd__nor4_1 _0954_ (.A(\cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[1] ),
    .Y(gfpga_pad_GPIO_PAD[9]));
 sky130_fd_sc_hd__nor4_1 _0955_ (.A(\cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_right_2__1_.GPIO_DIR[0] ),
    .Y(gfpga_pad_GPIO_PAD[8]));
 sky130_fd_sc_hd__nor4_1 _0956_ (.A(\cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[7] ),
    .Y(gfpga_pad_GPIO_PAD[23]));
 sky130_fd_sc_hd__nor4_1 _0957_ (.A(\cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[6] ),
    .Y(gfpga_pad_GPIO_PAD[22]));
 sky130_fd_sc_hd__nor4_1 _0958_ (.A(\cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[5] ),
    .Y(gfpga_pad_GPIO_PAD[21]));
 sky130_fd_sc_hd__nor4_1 _0959_ (.A(\cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[4] ),
    .Y(gfpga_pad_GPIO_PAD[20]));
 sky130_fd_sc_hd__nor4_1 _0960_ (.A(\cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[3] ),
    .Y(gfpga_pad_GPIO_PAD[19]));
 sky130_fd_sc_hd__nor4_1 _0961_ (.A(\cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[2] ),
    .Y(gfpga_pad_GPIO_PAD[18]));
 sky130_fd_sc_hd__nor4_1 _0962_ (.A(\cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[1] ),
    .Y(gfpga_pad_GPIO_PAD[17]));
 sky130_fd_sc_hd__nor4_1 _0963_ (.A(\cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_bottom_1__0_.GPIO_DIR[0] ),
    .Y(gfpga_pad_GPIO_PAD[16]));
 sky130_fd_sc_hd__nor4_1 _0964_ (.A(\cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[7] ),
    .Y(gfpga_pad_GPIO_PAD[31]));
 sky130_fd_sc_hd__nor4_1 _0965_ (.A(\cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[6] ),
    .Y(gfpga_pad_GPIO_PAD[30]));
 sky130_fd_sc_hd__nor4_1 _0966_ (.A(\cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[5] ),
    .Y(gfpga_pad_GPIO_PAD[29]));
 sky130_fd_sc_hd__nor4_1 _0967_ (.A(\cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[4] ),
    .Y(gfpga_pad_GPIO_PAD[28]));
 sky130_fd_sc_hd__nor4_1 _0968_ (.A(\cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[3] ),
    .Y(gfpga_pad_GPIO_PAD[27]));
 sky130_fd_sc_hd__nor4_1 _0969_ (.A(\cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[2] ),
    .Y(gfpga_pad_GPIO_PAD[26]));
 sky130_fd_sc_hd__nor4_1 _0970_ (.A(\cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[1] ),
    .Y(gfpga_pad_GPIO_PAD[25]));
 sky130_fd_sc_hd__nor4_1 _0971_ (.A(\cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out ),
    .D(\grid_io_left_0__1_.GPIO_DIR[0] ),
    .Y(gfpga_pad_GPIO_PAD[24]));
 sky130_fd_sc_hd__nand2_1 _0972_ (.A(\sb_1__1_.Q_in[40] ),
    .B(\sb_1__1_.Q_in[41] ),
    .Y(_0528_));
 sky130_fd_sc_hd__or2_1 _0973_ (.A(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .B(_0528_),
    .X(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _0974_ (.A(\sb_0__1_.Q_in[66] ),
    .B(\sb_0__1_.Q_in[67] ),
    .Y(_0529_));
 sky130_fd_sc_hd__or3_1 _0975_ (.A(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .B(_0528_),
    .C(_0529_),
    .X(\cby_0__1_.mux_right_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _0976_ (.A(\sb_0__0_.Q_in[72] ),
    .B(\sb_0__0_.Q_in[73] ),
    .Y(_0530_));
 sky130_fd_sc_hd__or4_4 _0977_ (.A(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .B(_0528_),
    .C(_0529_),
    .D(_0530_),
    .X(\cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand3_1 _0978_ (.A(\sb_1__1_.Q_in[42] ),
    .B(\sb_1__1_.Q_in[43] ),
    .C(_0523_),
    .Y(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(\sb_0__1_.Q_in[64] ),
    .B(\sb_0__1_.Q_in[65] ),
    .Y(_0531_));
 sky130_fd_sc_hd__nor2_1 _0980_ (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .B(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_1 _0981_ (.A(_0532_),
    .Y(\cby_0__1_.mux_right_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand3_1 _0982_ (.A(\sb_0__0_.Q_in[70] ),
    .B(\sb_0__0_.Q_in[71] ),
    .C(_0532_),
    .Y(\cbx_1__0_.mux_top_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand2b_1 _0983_ (.A_N(\sb_1__0_.Q_in[13] ),
    .B(\sb_1__0_.Q_in[12] ),
    .Y(_0533_));
 sky130_fd_sc_hd__or2_1 _0984_ (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .B(_0533_),
    .X(\cby_1__1_.mux_left_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand2_1 _0985_ (.A(\sb_1__1_.Q_in[44] ),
    .B(\sb_1__1_.Q_in[45] ),
    .Y(_0534_));
 sky130_fd_sc_hd__or3_1 _0986_ (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .B(_0533_),
    .C(_0534_),
    .X(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(\sb_0__1_.Q_in[62] ),
    .B(\sb_0__1_.Q_in[63] ),
    .Y(_0535_));
 sky130_fd_sc_hd__nor4_4 _0988_ (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .B(_0533_),
    .C(_0534_),
    .D(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__inv_1 _0989_ (.A(_0536_),
    .Y(\cby_0__1_.mux_right_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand3_1 _0990_ (.A(\sb_0__0_.Q_in[68] ),
    .B(\sb_0__0_.Q_in[69] ),
    .C(_0536_),
    .Y(\cbx_1__0_.mux_top_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand3b_1 _0991_ (.A_N(\sb_1__0_.Q_in[78] ),
    .B(\sb_1__0_.Q_in[79] ),
    .C(_0526_),
    .Y(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__or3b_1 _0992_ (.A(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_5_.out ),
    .B(\sb_0__0_.Q_in[30] ),
    .C_N(\sb_0__0_.Q_in[31] ),
    .X(\cby_0__1_.mux_right_ipin_3.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand3_1 _0993_ (.A(\sb_0__1_.Q_in[68] ),
    .B(\sb_0__1_.Q_in[69] ),
    .C(_0525_),
    .Y(\cby_0__1_.mux_right_ipin_3.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _0994_ (.A(\sb_0__0_.Q_in[74] ),
    .B(\cby_0__1_.mux_right_ipin_3.INVTX1_5_.out ),
    .Y(_0537_));
 sky130_fd_sc_hd__o211ai_1 _0995_ (.A1(\sb_0__0_.Q_in[74] ),
    .A2(_0526_),
    .B1(_0537_),
    .C1(\sb_0__0_.Q_in[75] ),
    .Y(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand3_1 _0996_ (.A(\sb_0__0_.Q_in[66] ),
    .B(\sb_0__0_.Q_in[67] ),
    .C(_0520_),
    .Y(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand2b_1 _0997_ (.A_N(\sb_1__0_.Q_in[21] ),
    .B(\sb_1__0_.Q_in[20] ),
    .Y(_0538_));
 sky130_fd_sc_hd__nor2_1 _0998_ (.A(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.out ),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__inv_1 _0999_ (.A(_0539_),
    .Y(\cby_1__1_.mux_left_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand3_1 _1000_ (.A(\sb_1__1_.Q_in[56] ),
    .B(\sb_1__1_.Q_in[57] ),
    .C(_0539_),
    .Y(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1001_ (.A(\sb_1__1_.Q_in[56] ),
    .B(\sb_1__1_.Q_in[57] ),
    .Y(_0540_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(\sb_0__1_.Q_in[50] ),
    .B(\sb_0__1_.Q_in[51] ),
    .Y(_0541_));
 sky130_fd_sc_hd__nor4_1 _1003_ (.A(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.out ),
    .B(_0538_),
    .C(_0540_),
    .D(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_1 _1004_ (.A(_0542_),
    .Y(\cby_0__1_.mux_right_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__and2_0 _1005_ (.A(\sb_0__0_.Q_in[52] ),
    .B(\sb_0__0_.Q_in[53] ),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _1006_ (.A(_0542_),
    .B(_0543_),
    .Y(\cbx_1__0_.mux_top_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand2_1 _1007_ (.A(\sb_1__1_.Q_in[59] ),
    .B(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.out ),
    .Y(_0544_));
 sky130_fd_sc_hd__o211ai_1 _1008_ (.A1(\sb_1__1_.Q_in[59] ),
    .A2(_0527_),
    .B1(_0544_),
    .C1(\sb_1__1_.Q_in[58] ),
    .Y(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1009_ (.A(\sb_0__1_.Q_in[48] ),
    .B(\sb_0__1_.Q_in[49] ),
    .Y(_0545_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .B(_0545_),
    .X(\cby_0__1_.mux_right_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _1011_ (.A(\sb_0__0_.Q_in[50] ),
    .B(\sb_0__0_.Q_in[51] ),
    .Y(_0546_));
 sky130_fd_sc_hd__or3_1 _1012_ (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .B(_0545_),
    .C(_0546_),
    .X(\cbx_1__0_.mux_top_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__nor2b_1 _1013_ (.A(\sb_1__0_.Q_in[29] ),
    .B_N(\sb_1__0_.Q_in[28] ),
    .Y(_0547_));
 sky130_fd_sc_hd__nand3_1 _1014_ (.A(_0542_),
    .B(_0543_),
    .C(_0547_),
    .Y(\cby_1__1_.mux_left_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__and2_0 _1015_ (.A(\sb_1__1_.Q_in[60] ),
    .B(\sb_1__1_.Q_in[61] ),
    .X(_0548_));
 sky130_fd_sc_hd__nand4_1 _1016_ (.A(_0542_),
    .B(_0543_),
    .C(_0547_),
    .D(_0548_),
    .Y(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1017_ (.A(\sb_0__1_.Q_in[46] ),
    .B(\sb_0__1_.Q_in[47] ),
    .Y(_0549_));
 sky130_fd_sc_hd__or2_1 _1018_ (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_5_.out ),
    .B(_0549_),
    .X(\cby_0__1_.mux_right_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _1019_ (.A(\sb_0__0_.Q_in[48] ),
    .B(\sb_0__0_.Q_in[49] ),
    .Y(_0550_));
 sky130_fd_sc_hd__nor3_1 _1020_ (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_5_.out ),
    .B(_0549_),
    .C(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__inv_1 _1021_ (.A(_0551_),
    .Y(\cbx_1__0_.mux_top_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand3_1 _1022_ (.A(\sb_0__0_.Q_in[46] ),
    .B(\sb_0__0_.Q_in[47] ),
    .C(_0521_),
    .Y(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__nor2b_1 _1023_ (.A(\sb_0__0_.Q_in[33] ),
    .B_N(\sb_0__0_.Q_in[32] ),
    .Y(_0552_));
 sky130_fd_sc_hd__nand2_1 _1024_ (.A(_0522_),
    .B(_0552_),
    .Y(\cby_0__1_.mux_left_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__or3b_1 _1025_ (.A(\sb_0__1_.Q_in[15] ),
    .B(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.out ),
    .C_N(\sb_0__1_.Q_in[14] ),
    .X(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_2_.out ));
 sky130_fd_sc_hd__or3b_1 _1026_ (.A(\sb_1__1_.Q_in[13] ),
    .B(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_2_.out ),
    .C_N(\sb_1__1_.Q_in[12] ),
    .X(\cby_1__1_.mux_left_ipin_4.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _1027_ (.A(\sb_1__0_.Q_in[72] ),
    .B(\sb_1__0_.Q_in[73] ),
    .Y(_0553_));
 sky130_fd_sc_hd__or2_1 _1028_ (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_3_.out ),
    .B(_0553_),
    .X(\cbx_1__0_.mux_top_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__inv_1 _1029_ (.A(\sb_0__0_.Q_in[25] ),
    .Y(_0554_));
 sky130_fd_sc_hd__nor2_1 _1030_ (.A(_0554_),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .Y(_0555_));
 sky130_fd_sc_hd__o21ai_1 _1031_ (.A1(\sb_0__0_.Q_in[25] ),
    .A2(\cbx_1__0_.mux_top_ipin_0.INVTX1_5_.out ),
    .B1(\sb_0__0_.Q_in[24] ),
    .Y(_0556_));
 sky130_fd_sc_hd__o21ai_1 _1032_ (.A1(\sb_0__0_.Q_in[24] ),
    .A2(_0555_),
    .B1(_0556_),
    .Y(\cby_0__1_.mux_right_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__nor3b_1 _1033_ (.A(\sb_1__1_.Q_in[15] ),
    .B(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.out ),
    .C_N(\sb_1__1_.Q_in[14] ),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_1 _1034_ (.A(_0557_),
    .Y(\cby_1__1_.mux_left_ipin_5.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand3_1 _1035_ (.A(\sb_1__0_.Q_in[70] ),
    .B(\sb_1__0_.Q_in[71] ),
    .C(_0557_),
    .Y(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__or3b_1 _1036_ (.A(\sb_0__0_.Q_in[23] ),
    .B(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .C_N(\sb_0__0_.Q_in[22] ),
    .X(\cby_0__1_.mux_left_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__or3b_2 _1037_ (.A(\sb_0__0_.Q_in[15] ),
    .B(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.out ),
    .C_N(\sb_0__0_.Q_in[14] ),
    .X(\cby_0__1_.mux_right_ipin_3.INVTX1_2_.out ));
 sky130_fd_sc_hd__or4b_1 _1038_ (.A(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.out ),
    .C(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ),
    .D_N(\sb_0__1_.Q_in[31] ),
    .X(_0558_));
 sky130_fd_sc_hd__or2_1 _1039_ (.A(\sb_0__1_.Q_in[30] ),
    .B(_0558_),
    .X(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_4_.out ));
 sky130_fd_sc_hd__nor4b_2 _1040_ (.A(\sb_0__1_.Q_in[30] ),
    .B(_0558_),
    .C(\sb_1__1_.Q_in[28] ),
    .D_N(\sb_1__1_.Q_in[29] ),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_1 _1041_ (.A(_0559_),
    .Y(\cby_1__1_.mux_left_ipin_4.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand3_1 _1042_ (.A(\sb_1__0_.Q_in[52] ),
    .B(\sb_1__0_.Q_in[53] ),
    .C(_0559_),
    .Y(\cbx_1__0_.mux_top_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__nor2b_1 _1043_ (.A(\sb_0__0_.Q_in[9] ),
    .B_N(\sb_0__0_.Q_in[8] ),
    .Y(_0560_));
 sky130_fd_sc_hd__nand4_1 _1044_ (.A(\sb_1__0_.Q_in[52] ),
    .B(\sb_1__0_.Q_in[53] ),
    .C(_0559_),
    .D(_0560_),
    .Y(\cby_0__1_.mux_right_ipin_0.INVTX1_2_.out ));
 sky130_fd_sc_hd__or3b_1 _1045_ (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_2_.out ),
    .B(\sb_0__1_.Q_in[26] ),
    .C_N(\sb_0__1_.Q_in[27] ),
    .X(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand2b_1 _1046_ (.A_N(\sb_1__1_.Q_in[24] ),
    .B(\sb_1__1_.Q_in[25] ),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2b_1 _1047_ (.A_N(\sb_1__1_.Q_in[25] ),
    .B(\sb_1__1_.Q_in[24] ),
    .Y(_0562_));
 sky130_fd_sc_hd__o22ai_2 _1048_ (.A1(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .A2(_0561_),
    .B1(_0562_),
    .B2(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_4_.out ),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_1 _1049_ (.A(_0563_),
    .Y(\cby_1__1_.mux_left_ipin_2.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand3_1 _1050_ (.A(\sb_1__0_.Q_in[56] ),
    .B(\sb_1__0_.Q_in[57] ),
    .C(_0563_),
    .Y(\cbx_1__0_.mux_top_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__nor2b_1 _1051_ (.A(\sb_0__0_.Q_in[13] ),
    .B_N(\sb_0__0_.Q_in[12] ),
    .Y(_0564_));
 sky130_fd_sc_hd__nand4_1 _1052_ (.A(\sb_1__0_.Q_in[56] ),
    .B(\sb_1__0_.Q_in[57] ),
    .C(_0563_),
    .D(_0564_),
    .Y(\cby_0__1_.mux_right_ipin_2.INVTX1_2_.out ));
 sky130_fd_sc_hd__nor2b_1 _1053_ (.A(\sb_0__1_.Q_in[33] ),
    .B_N(\sb_0__1_.Q_in[32] ),
    .Y(_0565_));
 sky130_fd_sc_hd__nand3_1 _1054_ (.A(_0522_),
    .B(_0552_),
    .C(_0565_),
    .Y(\cbx_1__1_.mux_bottom_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__nor2b_1 _1055_ (.A(\sb_1__1_.Q_in[30] ),
    .B_N(\sb_1__1_.Q_in[31] ),
    .Y(_0566_));
 sky130_fd_sc_hd__nand4_1 _1056_ (.A(_0522_),
    .B(_0552_),
    .C(_0565_),
    .D(_0566_),
    .Y(\cby_1__1_.mux_left_ipin_5.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1057_ (.A(\sb_1__0_.Q_in[50] ),
    .B(\sb_1__0_.Q_in[51] ),
    .Y(_0567_));
 sky130_fd_sc_hd__or2_1 _1058_ (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_5_.out ),
    .B(_0567_),
    .X(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2b_1 _1059_ (.A_N(\sb_0__0_.Q_in[7] ),
    .B(\sb_0__0_.Q_in[6] ),
    .Y(_0568_));
 sky130_fd_sc_hd__or3_1 _1060_ (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_5_.out ),
    .B(_0567_),
    .C(_0568_),
    .X(\cby_0__1_.mux_left_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand2b_1 _1061_ (.A_N(\sb_0__1_.Q_in[28] ),
    .B(\sb_0__1_.Q_in[29] ),
    .Y(_0569_));
 sky130_fd_sc_hd__nor4_1 _1062_ (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_5_.out ),
    .B(_0567_),
    .C(_0568_),
    .D(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__inv_1 _1063_ (.A(_0570_),
    .Y(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_4_.out ));
 sky130_fd_sc_hd__nor2b_1 _1064_ (.A(\sb_1__1_.Q_in[26] ),
    .B_N(\sb_1__1_.Q_in[27] ),
    .Y(_0571_));
 sky130_fd_sc_hd__nand2_1 _1065_ (.A(_0570_),
    .B(_0571_),
    .Y(\cby_1__1_.mux_left_ipin_3.INVTX1_5_.out ));
 sky130_fd_sc_hd__and2_0 _1066_ (.A(\sb_1__0_.Q_in[54] ),
    .B(\sb_1__0_.Q_in[55] ),
    .X(_0572_));
 sky130_fd_sc_hd__nand3_1 _1067_ (.A(_0570_),
    .B(_0571_),
    .C(_0572_),
    .Y(\cbx_1__0_.mux_top_ipin_1.INVTX1_3_.out ));
 sky130_fd_sc_hd__nor2b_1 _1068_ (.A(\sb_0__0_.Q_in[11] ),
    .B_N(\sb_0__0_.Q_in[10] ),
    .Y(_0573_));
 sky130_fd_sc_hd__nand4_1 _1069_ (.A(_0570_),
    .B(_0571_),
    .C(_0572_),
    .D(_0573_),
    .Y(\cby_0__1_.mux_right_ipin_1.INVTX1_2_.out ));
 sky130_fd_sc_hd__nor3b_1 _1070_ (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .B(\sb_1__0_.Q_in[34] ),
    .C_N(\sb_1__0_.Q_in[35] ),
    .Y(_0574_));
 sky130_fd_sc_hd__inv_1 _1071_ (.A(_0574_),
    .Y(\cby_1__1_.mux_left_ipin_5.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand3_1 _1072_ (.A(\sb_1__1_.Q_in[66] ),
    .B(\sb_1__1_.Q_in[67] ),
    .C(_0574_),
    .Y(\cbx_1__1_.mux_bottom_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1073_ (.A(\sb_0__1_.Q_in[70] ),
    .B(\sb_0__1_.Q_in[71] ),
    .Y(_0575_));
 sky130_fd_sc_hd__or2_1 _1074_ (.A(\cbx_1__1_.mux_bottom_ipin_0.INVTX1_5_.out ),
    .B(_0575_),
    .X(\cby_0__1_.mux_left_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__nor2b_1 _1075_ (.A(\sb_1__0_.Q_in[17] ),
    .B_N(\sb_1__0_.Q_in[16] ),
    .Y(_0576_));
 sky130_fd_sc_hd__and4_1 _1076_ (.A(\sb_0__0_.Q_in[68] ),
    .B(\sb_0__0_.Q_in[69] ),
    .C(_0536_),
    .D(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__inv_1 _1077_ (.A(_0577_),
    .Y(\cby_1__1_.mux_left_ipin_4.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand3_2 _1078_ (.A(\sb_1__1_.Q_in[48] ),
    .B(\sb_1__1_.Q_in[49] ),
    .C(_0577_),
    .Y(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _1079_ (.A(\sb_0__1_.Q_in[54] ),
    .B(\sb_0__1_.Q_in[55] ),
    .Y(_0578_));
 sky130_fd_sc_hd__or2_1 _1080_ (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_3_.out ),
    .B(_0578_),
    .X(\cby_0__1_.mux_left_ipin_0.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand3_1 _1081_ (.A(\sb_0__1_.Q_in[52] ),
    .B(\sb_0__1_.Q_in[53] ),
    .C(_0524_),
    .Y(\cby_0__1_.mux_right_ipin_3.INVTX1_3_.out ));
 sky130_fd_sc_hd__nand2_1 _1082_ (.A(\sb_0__1_.Q_in[25] ),
    .B(_0527_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2b_1 _1083_ (.A_N(\sb_0__1_.Q_in[25] ),
    .B(\sb_0__1_.Q_in[24] ),
    .Y(_0580_));
 sky130_fd_sc_hd__o22a_1 _1084_ (.A1(\sb_0__1_.Q_in[24] ),
    .A2(_0579_),
    .B1(_0580_),
    .B2(\cby_0__1_.mux_right_ipin_1.INVTX1_2_.out ),
    .X(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand2_1 _1085_ (.A(\sb_1__0_.Q_in[56] ),
    .B(\sb_1__0_.Q_in[57] ),
    .Y(_0581_));
 sky130_fd_sc_hd__nor2b_1 _1086_ (.A(\sb_0__1_.Q_in[23] ),
    .B_N(\sb_0__1_.Q_in[22] ),
    .Y(_0582_));
 sky130_fd_sc_hd__nand4b_1 _1087_ (.A_N(_0581_),
    .B(_0564_),
    .C(_0582_),
    .D(_0563_),
    .Y(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_4_.out ));
 sky130_fd_sc_hd__or3b_2 _1088_ (.A(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.out ),
    .B(\sb_1__0_.Q_in[36] ),
    .C_N(\sb_1__0_.Q_in[37] ),
    .X(\cby_1__1_.mux_left_ipin_0.INVTX1_4_.out ));
 sky130_fd_sc_hd__nand3b_1 _1089_ (.A_N(\sb_1__0_.Q_in[32] ),
    .B(\sb_1__0_.Q_in[33] ),
    .C(_0551_),
    .Y(\cby_1__1_.mux_left_ipin_4.INVTX1_4_.out ));
 sky130_fd_sc_hd__or3b_1 _1090_ (.A(\cbx_1__0_.mux_top_ipin_1.INVTX1_2_.out ),
    .B(\sb_1__0_.Q_in[30] ),
    .C_N(\sb_1__0_.Q_in[31] ),
    .X(\cby_1__1_.mux_left_ipin_3.INVTX1_4_.out ));
 sky130_fd_sc_hd__or3b_1 _1091_ (.A(\sb_1__0_.Q_in[19] ),
    .B(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .C_N(\sb_1__0_.Q_in[18] ),
    .X(\cby_1__1_.mux_left_ipin_5.INVTX1_2_.out ));
 sky130_fd_sc_hd__or3b_1 _1092_ (.A(\sb_1__0_.Q_in[15] ),
    .B(\cbx_1__0_.mux_top_ipin_1.INVTX1_4_.out ),
    .C_N(\sb_1__0_.Q_in[14] ),
    .X(\cby_1__1_.mux_left_ipin_3.INVTX1_2_.out ));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(\sb_1__1_.Q_in[64] ),
    .B(\sb_1__1_.Q_in[65] ),
    .Y(_0583_));
 sky130_fd_sc_hd__or2_1 _1094_ (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_4_.out ),
    .B(_0583_),
    .X(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1095_ (.A(\sb_1__1_.Q_in[62] ),
    .B(\sb_1__1_.Q_in[63] ),
    .Y(_0584_));
 sky130_fd_sc_hd__or2_1 _1096_ (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_4_.out ),
    .B(_0584_),
    .X(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1097_ (.A(\sb_1__1_.Q_in[46] ),
    .B(\sb_1__1_.Q_in[47] ),
    .Y(_0585_));
 sky130_fd_sc_hd__or2_1 _1098_ (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_2_.out ),
    .B(_0585_),
    .X(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_3_.out ));
 sky130_fd_sc_hd__or3b_2 _1099_ (.A(\sb_1__1_.Q_in[33] ),
    .B(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.out ),
    .C_N(\sb_1__1_.Q_in[32] ),
    .X(\cby_1__1_.mux_left_ipin_0.INVTX1_5_.out ));
 sky130_fd_sc_hd__or3b_1 _1100_ (.A(\sb_1__1_.Q_in[23] ),
    .B(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .C_N(\sb_1__1_.Q_in[22] ),
    .X(\cby_1__1_.mux_left_ipin_1.INVTX1_5_.out ));
 sky130_fd_sc_hd__nand2_1 _1103_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2b_1 _1104_ (.A_N(wl_address[0]),
    .B(enable),
    .Y(_0589_));
 sky130_fd_sc_hd__or3b_2 _1107_ (.A(_0589_),
    .B(wl_address[1]),
    .C_N(wl_address[2]),
    .X(_0592_));
 sky130_fd_sc_hd__nor2_1 _1108_ (.A(_0588_),
    .B(_0592_),
    .Y(\cbx_1__0_.wl[38] ));
 sky130_fd_sc_hd__nand2b_1 _1109_ (.A_N(wl_address[2]),
    .B(wl_address[1]),
    .Y(_0593_));
 sky130_fd_sc_hd__nand2_1 _1111_ (.A(wl_address[0]),
    .B(enable),
    .Y(_0595_));
 sky130_fd_sc_hd__nor3_1 _1113_ (.A(_0588_),
    .B(_0593_),
    .C(_0595_),
    .Y(\cbx_1__0_.wl[37] ));
 sky130_fd_sc_hd__nor3_1 _1115_ (.A(_0588_),
    .B(_0589_),
    .C(_0593_),
    .Y(\cbx_1__0_.wl[36] ));
 sky130_fd_sc_hd__nor4_1 _1116_ (.A(wl_address[1]),
    .B(wl_address[2]),
    .C(_0588_),
    .D(_0595_),
    .Y(\cbx_1__0_.wl[35] ));
 sky130_fd_sc_hd__nor4_1 _1117_ (.A(wl_address[1]),
    .B(wl_address[2]),
    .C(_0588_),
    .D(_0589_),
    .Y(\cbx_1__0_.wl[34] ));
 sky130_fd_sc_hd__nand2_1 _1118_ (.A(wl_address[1]),
    .B(wl_address[2]),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2b_1 _1119_ (.A_N(wl_address[3]),
    .B(wl_address[4]),
    .Y(_0599_));
 sky130_fd_sc_hd__nor3_1 _1121_ (.A(_0595_),
    .B(_0598_),
    .C(_0599_),
    .Y(\cbx_1__0_.wl[33] ));
 sky130_fd_sc_hd__nor3_1 _1122_ (.A(_0589_),
    .B(_0598_),
    .C(_0599_),
    .Y(\cbx_1__0_.wl[32] ));
 sky130_fd_sc_hd__nand4b_1 _1123_ (.A_N(wl_address[1]),
    .B(wl_address[2]),
    .C(wl_address[0]),
    .D(enable),
    .Y(_0601_));
 sky130_fd_sc_hd__nor2_1 _1124_ (.A(_0599_),
    .B(_0601_),
    .Y(\cbx_1__0_.wl[2] ));
 sky130_fd_sc_hd__nor2_1 _1125_ (.A(_0592_),
    .B(_0599_),
    .Y(\cbx_1__0_.wl[1] ));
 sky130_fd_sc_hd__nor3_1 _1126_ (.A(_0593_),
    .B(_0595_),
    .C(_0599_),
    .Y(\cbx_1__0_.wl[0] ));
 sky130_fd_sc_hd__nor3_1 _1127_ (.A(_0589_),
    .B(_0593_),
    .C(_0599_),
    .Y(\cbx_1__0_.wl[28] ));
 sky130_fd_sc_hd__nor4_1 _1128_ (.A(wl_address[1]),
    .B(wl_address[2]),
    .C(_0595_),
    .D(_0599_),
    .Y(\cbx_1__0_.wl[27] ));
 sky130_fd_sc_hd__nor4_1 _1129_ (.A(wl_address[1]),
    .B(wl_address[2]),
    .C(_0589_),
    .D(_0599_),
    .Y(\cbx_1__0_.wl[26] ));
 sky130_fd_sc_hd__nand2b_1 _1130_ (.A_N(wl_address[4]),
    .B(wl_address[3]),
    .Y(_0602_));
 sky130_fd_sc_hd__nor3_1 _1132_ (.A(_0595_),
    .B(_0598_),
    .C(_0602_),
    .Y(\cbx_1__0_.wl[25] ));
 sky130_fd_sc_hd__nor3_1 _1133_ (.A(_0589_),
    .B(_0598_),
    .C(_0602_),
    .Y(\cbx_1__0_.wl[24] ));
 sky130_fd_sc_hd__nor2_1 _1134_ (.A(_0601_),
    .B(_0602_),
    .Y(\cbx_1__0_.wl[23] ));
 sky130_fd_sc_hd__nor2_1 _1135_ (.A(_0592_),
    .B(_0602_),
    .Y(\cbx_1__0_.wl[22] ));
 sky130_fd_sc_hd__nor3_1 _1136_ (.A(_0593_),
    .B(_0595_),
    .C(_0602_),
    .Y(\cbx_1__0_.wl[21] ));
 sky130_fd_sc_hd__nor3_1 _1137_ (.A(_0589_),
    .B(_0593_),
    .C(_0602_),
    .Y(\cbx_1__0_.wl[20] ));
 sky130_fd_sc_hd__nor4_1 _1138_ (.A(wl_address[1]),
    .B(wl_address[2]),
    .C(_0595_),
    .D(_0602_),
    .Y(\cbx_1__0_.wl[19] ));
 sky130_fd_sc_hd__nor4_1 _1139_ (.A(wl_address[1]),
    .B(wl_address[2]),
    .C(_0589_),
    .D(_0602_),
    .Y(\cbx_1__0_.wl[18] ));
 sky130_fd_sc_hd__nor4_1 _1140_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .C(_0595_),
    .D(_0598_),
    .Y(\cbx_1__0_.wl[17] ));
 sky130_fd_sc_hd__nor4_1 _1141_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .C(_0589_),
    .D(_0598_),
    .Y(\cbx_1__0_.wl[16] ));
 sky130_fd_sc_hd__nor3_1 _1142_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .C(_0601_),
    .Y(\cbx_1__0_.wl[15] ));
 sky130_fd_sc_hd__nor3_1 _1143_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .C(_0592_),
    .Y(\cbx_1__0_.wl[14] ));
 sky130_fd_sc_hd__nor4_1 _1144_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .C(_0593_),
    .D(_0595_),
    .Y(\cbx_1__0_.wl[13] ));
 sky130_fd_sc_hd__nor4_1 _1145_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .C(_0589_),
    .D(_0593_),
    .Y(\cbx_1__0_.wl[12] ));
 sky130_fd_sc_hd__or4_1 _1146_ (.A(wl_address[4]),
    .B(wl_address[3]),
    .C(wl_address[1]),
    .D(wl_address[2]),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _1147_ (.A(_0595_),
    .B(_0604_),
    .Y(\cbx_1__0_.wl[11] ));
 sky130_fd_sc_hd__nor2_1 _1148_ (.A(_0589_),
    .B(_0604_),
    .Y(\cbx_1__0_.wl[10] ));
 sky130_fd_sc_hd__or4_1 _1149_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0605_));
 sky130_fd_sc_hd__nand2_1 _1151_ (.A(\grid_clb_1__1_.Q_in[5] ),
    .B(_0605_),
    .Y(_0607_));
 sky130_fd_sc_hd__nor4_1 _1152_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _1153_ (.A(\grid_clb_1__1_.Q_in[1] ),
    .B(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor4_1 _1154_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0610_));
 sky130_fd_sc_hd__a21oi_1 _1155_ (.A1(_0607_),
    .A2(_0609_),
    .B1(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_1 _1156_ (.A(\grid_clb_1__1_.Q_in[4] ),
    .B(_0608_),
    .Y(_0612_));
 sky130_fd_sc_hd__o21ai_1 _1157_ (.A1(\grid_clb_1__1_.Q_in[0] ),
    .A2(_0605_),
    .B1(_0610_),
    .Y(_0613_));
 sky130_fd_sc_hd__nor4_1 _1158_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0614_));
 sky130_fd_sc_hd__o21ai_0 _1159_ (.A1(_0612_),
    .A2(_0613_),
    .B1(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__nor2_1 _1160_ (.A(_0611_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__nand2_1 _1161_ (.A(\grid_clb_1__1_.Q_in[13] ),
    .B(_0605_),
    .Y(_0617_));
 sky130_fd_sc_hd__a21oi_1 _1162_ (.A1(\grid_clb_1__1_.Q_in[9] ),
    .A2(_0608_),
    .B1(_0610_),
    .Y(_0618_));
 sky130_fd_sc_hd__nand2_1 _1163_ (.A(\grid_clb_1__1_.Q_in[8] ),
    .B(_0608_),
    .Y(_0619_));
 sky130_fd_sc_hd__or4_1 _1164_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0620_));
 sky130_fd_sc_hd__a21oi_1 _1165_ (.A1(\grid_clb_1__1_.Q_in[12] ),
    .A2(_0605_),
    .B1(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__a22oi_1 _1166_ (.A1(_0617_),
    .A2(_0618_),
    .B1(_0619_),
    .B2(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nor4_1 _1167_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0623_));
 sky130_fd_sc_hd__o21ai_0 _1168_ (.A1(_0614_),
    .A2(_0622_),
    .B1(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _1169_ (.A(\grid_clb_1__1_.Q_in[11] ),
    .B(_0608_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand2_1 _1170_ (.A(\grid_clb_1__1_.Q_in[15] ),
    .B(_0605_),
    .Y(_0626_));
 sky130_fd_sc_hd__nand2_1 _1171_ (.A(\grid_clb_1__1_.Q_in[10] ),
    .B(_0608_),
    .Y(_0627_));
 sky130_fd_sc_hd__a21oi_1 _1172_ (.A1(\grid_clb_1__1_.Q_in[14] ),
    .A2(_0605_),
    .B1(_0620_),
    .Y(_0628_));
 sky130_fd_sc_hd__a32oi_1 _1173_ (.A1(_0620_),
    .A2(_0625_),
    .A3(_0626_),
    .B1(_0627_),
    .B2(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__mux2i_1 _1174_ (.A0(\grid_clb_1__1_.Q_in[3] ),
    .A1(\grid_clb_1__1_.Q_in[7] ),
    .S(_0605_),
    .Y(_0630_));
 sky130_fd_sc_hd__o21ai_0 _1175_ (.A1(\grid_clb_1__1_.Q_in[2] ),
    .A2(_0605_),
    .B1(_0610_),
    .Y(_0631_));
 sky130_fd_sc_hd__nor2_1 _1176_ (.A(\grid_clb_1__1_.Q_in[6] ),
    .B(_0608_),
    .Y(_0632_));
 sky130_fd_sc_hd__o221ai_1 _1177_ (.A1(_0610_),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0632_),
    .C1(_0614_),
    .Y(_0633_));
 sky130_fd_sc_hd__o21ai_0 _1178_ (.A1(_0614_),
    .A2(_0629_),
    .B1(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__o22a_1 _1179_ (.A1(_0616_),
    .A2(_0624_),
    .B1(_0634_),
    .B2(_0623_),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__inv_1 _1180_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_ff_0.DFFSRQ_0_.D ));
 sky130_fd_sc_hd__or4_1 _1181_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0635_));
 sky130_fd_sc_hd__nor4_1 _1182_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0636_));
 sky130_fd_sc_hd__nor4_1 _1183_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0637_));
 sky130_fd_sc_hd__nor2_1 _1184_ (.A(\grid_clb_1__1_.Q_in[32] ),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__or4_1 _1185_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0639_));
 sky130_fd_sc_hd__nor2_1 _1187_ (.A(\grid_clb_1__1_.Q_in[28] ),
    .B(_0639_),
    .Y(_0641_));
 sky130_fd_sc_hd__nor3_1 _1188_ (.A(_0636_),
    .B(_0638_),
    .C(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nor2_1 _1189_ (.A(\grid_clb_1__1_.Q_in[27] ),
    .B(_0639_),
    .Y(_0643_));
 sky130_fd_sc_hd__o21ai_0 _1190_ (.A1(\grid_clb_1__1_.Q_in[31] ),
    .A2(_0637_),
    .B1(_0636_),
    .Y(_0644_));
 sky130_fd_sc_hd__nor2_1 _1191_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__nand2_1 _1192_ (.A(\grid_clb_1__1_.Q_in[30] ),
    .B(_0637_),
    .Y(_0646_));
 sky130_fd_sc_hd__nand2_1 _1193_ (.A(\grid_clb_1__1_.Q_in[34] ),
    .B(_0639_),
    .Y(_0647_));
 sky130_fd_sc_hd__a21oi_1 _1194_ (.A1(_0646_),
    .A2(_0647_),
    .B1(_0636_),
    .Y(_0648_));
 sky130_fd_sc_hd__nor2_1 _1195_ (.A(\grid_clb_1__1_.Q_in[33] ),
    .B(_0637_),
    .Y(_0649_));
 sky130_fd_sc_hd__o21ai_0 _1196_ (.A1(\grid_clb_1__1_.Q_in[29] ),
    .A2(_0639_),
    .B1(_0636_),
    .Y(_0650_));
 sky130_fd_sc_hd__o21ai_0 _1197_ (.A1(_0649_),
    .A2(_0650_),
    .B1(_0635_),
    .Y(_0651_));
 sky130_fd_sc_hd__o32ai_1 _1198_ (.A1(_0635_),
    .A2(_0642_),
    .A3(_0645_),
    .B1(_0648_),
    .B2(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__nand2_1 _1199_ (.A(\grid_clb_1__1_.Q_in[19] ),
    .B(_0637_),
    .Y(_0653_));
 sky130_fd_sc_hd__nand2_1 _1200_ (.A(\grid_clb_1__1_.Q_in[23] ),
    .B(_0639_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_1 _1201_ (.A(\grid_clb_1__1_.Q_in[24] ),
    .B(_0639_),
    .Y(_0655_));
 sky130_fd_sc_hd__a21oi_1 _1202_ (.A1(\grid_clb_1__1_.Q_in[20] ),
    .A2(_0637_),
    .B1(_0636_),
    .Y(_0656_));
 sky130_fd_sc_hd__a32oi_1 _1203_ (.A1(_0636_),
    .A2(_0653_),
    .A3(_0654_),
    .B1(_0655_),
    .B2(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _1204_ (.A(\grid_clb_1__1_.Q_in[21] ),
    .B(_0637_),
    .Y(_0658_));
 sky130_fd_sc_hd__nand2_1 _1205_ (.A(\grid_clb_1__1_.Q_in[25] ),
    .B(_0639_),
    .Y(_0659_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(\grid_clb_1__1_.Q_in[22] ),
    .B(_0637_),
    .Y(_0660_));
 sky130_fd_sc_hd__a21oi_1 _1207_ (.A1(\grid_clb_1__1_.Q_in[26] ),
    .A2(_0639_),
    .B1(_0636_),
    .Y(_0661_));
 sky130_fd_sc_hd__a32oi_1 _1208_ (.A1(_0636_),
    .A2(_0658_),
    .A3(_0659_),
    .B1(_0660_),
    .B2(_0661_),
    .Y(_0662_));
 sky130_fd_sc_hd__mux2i_1 _1209_ (.A0(_0657_),
    .A1(_0662_),
    .S(_0635_),
    .Y(_0663_));
 sky130_fd_sc_hd__nor4_1 _1210_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0664_));
 sky130_fd_sc_hd__mux2_2 _1211_ (.A0(_0652_),
    .A1(_0663_),
    .S(_0664_),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__inv_2 _1212_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_ff_0.DFFSRQ_0_.D ));
 sky130_fd_sc_hd__or4_1 _1213_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0665_));
 sky130_fd_sc_hd__nor4_1 _1214_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0666_));
 sky130_fd_sc_hd__nor4_1 _1215_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0667_));
 sky130_fd_sc_hd__nor2_1 _1216_ (.A(\grid_clb_1__1_.Q_in[51] ),
    .B(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__or4_1 _1217_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0669_));
 sky130_fd_sc_hd__nor2_1 _1219_ (.A(\grid_clb_1__1_.Q_in[47] ),
    .B(_0669_),
    .Y(_0671_));
 sky130_fd_sc_hd__nor3_1 _1220_ (.A(_0666_),
    .B(_0668_),
    .C(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__nor2_1 _1221_ (.A(\grid_clb_1__1_.Q_in[46] ),
    .B(_0669_),
    .Y(_0673_));
 sky130_fd_sc_hd__o21ai_0 _1222_ (.A1(\grid_clb_1__1_.Q_in[50] ),
    .A2(_0667_),
    .B1(_0666_),
    .Y(_0674_));
 sky130_fd_sc_hd__nor2_1 _1223_ (.A(_0673_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__nand2_1 _1224_ (.A(\grid_clb_1__1_.Q_in[49] ),
    .B(_0667_),
    .Y(_0676_));
 sky130_fd_sc_hd__nand2_1 _1225_ (.A(\grid_clb_1__1_.Q_in[53] ),
    .B(_0669_),
    .Y(_0677_));
 sky130_fd_sc_hd__a21oi_1 _1226_ (.A1(_0676_),
    .A2(_0677_),
    .B1(_0666_),
    .Y(_0678_));
 sky130_fd_sc_hd__nor2_1 _1227_ (.A(\grid_clb_1__1_.Q_in[52] ),
    .B(_0667_),
    .Y(_0679_));
 sky130_fd_sc_hd__o21ai_0 _1228_ (.A1(\grid_clb_1__1_.Q_in[48] ),
    .A2(_0669_),
    .B1(_0666_),
    .Y(_0680_));
 sky130_fd_sc_hd__o21ai_0 _1229_ (.A1(_0679_),
    .A2(_0680_),
    .B1(_0665_),
    .Y(_0681_));
 sky130_fd_sc_hd__o32ai_1 _1230_ (.A1(_0665_),
    .A2(_0672_),
    .A3(_0675_),
    .B1(_0678_),
    .B2(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__nand2_1 _1231_ (.A(\grid_clb_1__1_.Q_in[38] ),
    .B(_0667_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _1232_ (.A(\grid_clb_1__1_.Q_in[42] ),
    .B(_0669_),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _1233_ (.A(\grid_clb_1__1_.Q_in[43] ),
    .B(_0669_),
    .Y(_0685_));
 sky130_fd_sc_hd__a21oi_1 _1234_ (.A1(\grid_clb_1__1_.Q_in[39] ),
    .A2(_0667_),
    .B1(_0666_),
    .Y(_0686_));
 sky130_fd_sc_hd__a32oi_1 _1235_ (.A1(_0666_),
    .A2(_0683_),
    .A3(_0684_),
    .B1(_0685_),
    .B2(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(\grid_clb_1__1_.Q_in[40] ),
    .B(_0667_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2_1 _1237_ (.A(\grid_clb_1__1_.Q_in[44] ),
    .B(_0669_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _1238_ (.A(\grid_clb_1__1_.Q_in[41] ),
    .B(_0667_),
    .Y(_0690_));
 sky130_fd_sc_hd__a21oi_1 _1239_ (.A1(\grid_clb_1__1_.Q_in[45] ),
    .A2(_0669_),
    .B1(_0666_),
    .Y(_0691_));
 sky130_fd_sc_hd__a32oi_1 _1240_ (.A1(_0666_),
    .A2(_0688_),
    .A3(_0689_),
    .B1(_0690_),
    .B2(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__mux2i_1 _1241_ (.A0(_0687_),
    .A1(_0692_),
    .S(_0665_),
    .Y(_0693_));
 sky130_fd_sc_hd__nor4_1 _1242_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0694_));
 sky130_fd_sc_hd__mux2_2 _1243_ (.A0(_0682_),
    .A1(_0693_),
    .S(_0694_),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__inv_2 _1244_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_ff_0.DFFSRQ_0_.D ));
 sky130_fd_sc_hd__or4_1 _1245_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_1 _1247_ (.A(\grid_clb_1__1_.Q_in[62] ),
    .B(_0695_),
    .Y(_0697_));
 sky130_fd_sc_hd__nor4_1 _1248_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0698_));
 sky130_fd_sc_hd__nand2_1 _1249_ (.A(\grid_clb_1__1_.Q_in[58] ),
    .B(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__nor4_1 _1250_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0700_));
 sky130_fd_sc_hd__a21oi_1 _1251_ (.A1(_0697_),
    .A2(_0699_),
    .B1(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__nor2_1 _1252_ (.A(\grid_clb_1__1_.Q_in[61] ),
    .B(_0698_),
    .Y(_0702_));
 sky130_fd_sc_hd__o21ai_1 _1253_ (.A1(\grid_clb_1__1_.Q_in[57] ),
    .A2(_0695_),
    .B1(_0700_),
    .Y(_0703_));
 sky130_fd_sc_hd__nor4_1 _1254_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0704_));
 sky130_fd_sc_hd__o21ai_0 _1255_ (.A1(_0702_),
    .A2(_0703_),
    .B1(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__nor2_1 _1256_ (.A(_0701_),
    .B(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _1257_ (.A(\grid_clb_1__1_.Q_in[70] ),
    .B(_0695_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21oi_1 _1258_ (.A1(\grid_clb_1__1_.Q_in[66] ),
    .A2(_0698_),
    .B1(_0700_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _1259_ (.A(\grid_clb_1__1_.Q_in[65] ),
    .B(_0698_),
    .Y(_0709_));
 sky130_fd_sc_hd__or4_1 _1260_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.out ),
    .X(_0710_));
 sky130_fd_sc_hd__a21oi_1 _1261_ (.A1(\grid_clb_1__1_.Q_in[69] ),
    .A2(_0695_),
    .B1(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__a22oi_1 _1262_ (.A1(_0707_),
    .A2(_0708_),
    .B1(_0709_),
    .B2(_0711_),
    .Y(_0712_));
 sky130_fd_sc_hd__nor4_1 _1263_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.out ),
    .B(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out ),
    .C(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.out ),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.out ),
    .Y(_0713_));
 sky130_fd_sc_hd__o21ai_0 _1264_ (.A1(_0704_),
    .A2(_0712_),
    .B1(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand2_1 _1265_ (.A(\grid_clb_1__1_.Q_in[68] ),
    .B(_0698_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand2_1 _1266_ (.A(\grid_clb_1__1_.Q_in[72] ),
    .B(_0695_),
    .Y(_0716_));
 sky130_fd_sc_hd__nand2_1 _1267_ (.A(\grid_clb_1__1_.Q_in[67] ),
    .B(_0698_),
    .Y(_0717_));
 sky130_fd_sc_hd__a21oi_1 _1268_ (.A1(\grid_clb_1__1_.Q_in[71] ),
    .A2(_0695_),
    .B1(_0710_),
    .Y(_0718_));
 sky130_fd_sc_hd__a32oi_1 _1269_ (.A1(_0710_),
    .A2(_0715_),
    .A3(_0716_),
    .B1(_0717_),
    .B2(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__mux2i_1 _1270_ (.A0(\grid_clb_1__1_.Q_in[60] ),
    .A1(\grid_clb_1__1_.Q_in[64] ),
    .S(_0695_),
    .Y(_0720_));
 sky130_fd_sc_hd__o21ai_0 _1271_ (.A1(\grid_clb_1__1_.Q_in[59] ),
    .A2(_0695_),
    .B1(_0700_),
    .Y(_0721_));
 sky130_fd_sc_hd__nor2_1 _1272_ (.A(\grid_clb_1__1_.Q_in[63] ),
    .B(_0698_),
    .Y(_0722_));
 sky130_fd_sc_hd__o221ai_1 _1273_ (.A1(_0700_),
    .A2(_0720_),
    .B1(_0721_),
    .B2(_0722_),
    .C1(_0704_),
    .Y(_0723_));
 sky130_fd_sc_hd__o21ai_1 _1274_ (.A1(_0704_),
    .A2(_0719_),
    .B1(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__o22a_1 _1275_ (.A1(_0706_),
    .A2(_0714_),
    .B1(_0724_),
    .B2(_0713_),
    .X(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ));
 sky130_fd_sc_hd__inv_1 _1276_ (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .Y(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_ff_0.DFFSRQ_0_.D ));
 sky130_fd_sc_hd__inv_1 _1277_ (.A(\grid_clb_1__1_.Q_in[104] ),
    .Y(_0292_));
 sky130_fd_sc_hd__inv_1 _1278_ (.A(\grid_clb_1__1_.Q_in[105] ),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_1 _1279_ (.A(\grid_clb_1__1_.Q_in[106] ),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_1 _1280_ (.A(\grid_clb_1__1_.Q_in[107] ),
    .Y(_0295_));
 sky130_fd_sc_hd__inv_1 _1281_ (.A(\grid_clb_1__1_.Q_in[100] ),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_1 _1282_ (.A(\grid_clb_1__1_.Q_in[101] ),
    .Y(_0289_));
 sky130_fd_sc_hd__inv_1 _1283_ (.A(\grid_clb_1__1_.Q_in[102] ),
    .Y(_0290_));
 sky130_fd_sc_hd__inv_1 _1284_ (.A(\grid_clb_1__1_.Q_in[103] ),
    .Y(_0291_));
 sky130_fd_sc_hd__inv_1 _1285_ (.A(\grid_clb_1__1_.Q_in[112] ),
    .Y(_0300_));
 sky130_fd_sc_hd__inv_1 _1286_ (.A(\grid_clb_1__1_.Q_in[113] ),
    .Y(_0301_));
 sky130_fd_sc_hd__inv_1 _1287_ (.A(\grid_clb_1__1_.Q_in[114] ),
    .Y(_0302_));
 sky130_fd_sc_hd__inv_1 _1288_ (.A(\grid_clb_1__1_.Q_in[115] ),
    .Y(_0303_));
 sky130_fd_sc_hd__inv_1 _1289_ (.A(\grid_clb_1__1_.Q_in[108] ),
    .Y(_0296_));
 sky130_fd_sc_hd__inv_1 _1290_ (.A(\grid_clb_1__1_.Q_in[109] ),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_1 _1291_ (.A(\grid_clb_1__1_.Q_in[110] ),
    .Y(_0298_));
 sky130_fd_sc_hd__inv_1 _1292_ (.A(\grid_clb_1__1_.Q_in[111] ),
    .Y(_0299_));
 sky130_fd_sc_hd__inv_1 _1293_ (.A(\grid_clb_1__1_.Q_in[120] ),
    .Y(_0308_));
 sky130_fd_sc_hd__inv_1 _1294_ (.A(\grid_clb_1__1_.Q_in[121] ),
    .Y(_0309_));
 sky130_fd_sc_hd__inv_1 _1295_ (.A(\grid_clb_1__1_.Q_in[122] ),
    .Y(_0310_));
 sky130_fd_sc_hd__inv_1 _1296_ (.A(\grid_clb_1__1_.Q_in[123] ),
    .Y(_0311_));
 sky130_fd_sc_hd__inv_1 _1297_ (.A(\grid_clb_1__1_.Q_in[116] ),
    .Y(_0304_));
 sky130_fd_sc_hd__inv_1 _1298_ (.A(\grid_clb_1__1_.Q_in[117] ),
    .Y(_0305_));
 sky130_fd_sc_hd__inv_1 _1299_ (.A(\grid_clb_1__1_.Q_in[118] ),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_1 _1300_ (.A(\grid_clb_1__1_.Q_in[119] ),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_1 _1301_ (.A(\grid_clb_1__1_.Q_in[128] ),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_1 _1302_ (.A(\grid_clb_1__1_.Q_in[129] ),
    .Y(_0317_));
 sky130_fd_sc_hd__inv_1 _1303_ (.A(\grid_clb_1__1_.Q_in[130] ),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_1 _1304_ (.A(\grid_clb_1__1_.Q_in[131] ),
    .Y(_0319_));
 sky130_fd_sc_hd__inv_1 _1305_ (.A(\grid_clb_1__1_.Q_in[124] ),
    .Y(_0312_));
 sky130_fd_sc_hd__inv_1 _1306_ (.A(\grid_clb_1__1_.Q_in[125] ),
    .Y(_0313_));
 sky130_fd_sc_hd__inv_1 _1307_ (.A(\grid_clb_1__1_.Q_in[126] ),
    .Y(_0314_));
 sky130_fd_sc_hd__inv_1 _1308_ (.A(\grid_clb_1__1_.Q_in[127] ),
    .Y(_0315_));
 sky130_fd_sc_hd__inv_1 _1309_ (.A(\grid_clb_1__1_.Q_in[136] ),
    .Y(_0324_));
 sky130_fd_sc_hd__inv_1 _1310_ (.A(\grid_clb_1__1_.Q_in[137] ),
    .Y(_0325_));
 sky130_fd_sc_hd__inv_1 _1311_ (.A(\grid_clb_1__1_.Q_in[138] ),
    .Y(_0326_));
 sky130_fd_sc_hd__inv_1 _1312_ (.A(\grid_clb_1__1_.Q_in[139] ),
    .Y(_0327_));
 sky130_fd_sc_hd__inv_1 _1313_ (.A(\grid_clb_1__1_.Q_in[132] ),
    .Y(_0320_));
 sky130_fd_sc_hd__inv_1 _1314_ (.A(\grid_clb_1__1_.Q_in[133] ),
    .Y(_0321_));
 sky130_fd_sc_hd__inv_1 _1315_ (.A(\grid_clb_1__1_.Q_in[134] ),
    .Y(_0322_));
 sky130_fd_sc_hd__inv_1 _1316_ (.A(\grid_clb_1__1_.Q_in[135] ),
    .Y(_0323_));
 sky130_fd_sc_hd__inv_1 _1317_ (.A(\grid_clb_1__1_.Q_in[144] ),
    .Y(_0332_));
 sky130_fd_sc_hd__inv_1 _1318_ (.A(\grid_clb_1__1_.Q_in[145] ),
    .Y(_0333_));
 sky130_fd_sc_hd__inv_1 _1319_ (.A(\grid_clb_1__1_.Q_in[146] ),
    .Y(_0334_));
 sky130_fd_sc_hd__inv_1 _1320_ (.A(\grid_clb_1__1_.Q_in[147] ),
    .Y(_0335_));
 sky130_fd_sc_hd__inv_1 _1321_ (.A(\grid_clb_1__1_.Q_in[140] ),
    .Y(_0328_));
 sky130_fd_sc_hd__inv_1 _1322_ (.A(\grid_clb_1__1_.Q_in[141] ),
    .Y(_0329_));
 sky130_fd_sc_hd__inv_1 _1323_ (.A(\grid_clb_1__1_.Q_in[142] ),
    .Y(_0330_));
 sky130_fd_sc_hd__inv_1 _1324_ (.A(\grid_clb_1__1_.Q_in[143] ),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_1 _1325_ (.A(\grid_clb_1__1_.Q_in[152] ),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_1 _1326_ (.A(\grid_clb_1__1_.Q_in[153] ),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_1 _1327_ (.A(\grid_clb_1__1_.Q_in[154] ),
    .Y(_0342_));
 sky130_fd_sc_hd__inv_1 _1328_ (.A(\grid_clb_1__1_.Q_in[155] ),
    .Y(_0343_));
 sky130_fd_sc_hd__inv_1 _1329_ (.A(\grid_clb_1__1_.Q_in[148] ),
    .Y(_0336_));
 sky130_fd_sc_hd__inv_1 _1330_ (.A(\grid_clb_1__1_.Q_in[149] ),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_1 _1331_ (.A(\grid_clb_1__1_.Q_in[150] ),
    .Y(_0338_));
 sky130_fd_sc_hd__inv_1 _1332_ (.A(\grid_clb_1__1_.Q_in[151] ),
    .Y(_0339_));
 sky130_fd_sc_hd__inv_1 _1333_ (.A(\grid_clb_1__1_.Q_in[160] ),
    .Y(_0348_));
 sky130_fd_sc_hd__inv_1 _1334_ (.A(\grid_clb_1__1_.Q_in[161] ),
    .Y(_0349_));
 sky130_fd_sc_hd__inv_1 _1335_ (.A(\grid_clb_1__1_.Q_in[162] ),
    .Y(_0350_));
 sky130_fd_sc_hd__inv_1 _1336_ (.A(\grid_clb_1__1_.Q_in[163] ),
    .Y(_0351_));
 sky130_fd_sc_hd__inv_1 _1337_ (.A(\grid_clb_1__1_.Q_in[156] ),
    .Y(_0344_));
 sky130_fd_sc_hd__inv_1 _1338_ (.A(\grid_clb_1__1_.Q_in[157] ),
    .Y(_0345_));
 sky130_fd_sc_hd__inv_1 _1339_ (.A(\grid_clb_1__1_.Q_in[158] ),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_1 _1340_ (.A(\grid_clb_1__1_.Q_in[159] ),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_1 _1341_ (.A(\grid_clb_1__1_.Q_in[168] ),
    .Y(_0356_));
 sky130_fd_sc_hd__inv_1 _1342_ (.A(\grid_clb_1__1_.Q_in[169] ),
    .Y(_0357_));
 sky130_fd_sc_hd__inv_1 _1343_ (.A(\grid_clb_1__1_.Q_in[170] ),
    .Y(_0358_));
 sky130_fd_sc_hd__inv_1 _1344_ (.A(\grid_clb_1__1_.Q_in[171] ),
    .Y(_0359_));
 sky130_fd_sc_hd__inv_1 _1345_ (.A(\grid_clb_1__1_.Q_in[164] ),
    .Y(_0352_));
 sky130_fd_sc_hd__inv_1 _1346_ (.A(\grid_clb_1__1_.Q_in[165] ),
    .Y(_0353_));
 sky130_fd_sc_hd__inv_1 _1347_ (.A(\grid_clb_1__1_.Q_in[166] ),
    .Y(_0354_));
 sky130_fd_sc_hd__inv_1 _1348_ (.A(\grid_clb_1__1_.Q_in[167] ),
    .Y(_0355_));
 sky130_fd_sc_hd__inv_1 _1349_ (.A(\grid_clb_1__1_.Q_in[176] ),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_1 _1350_ (.A(\grid_clb_1__1_.Q_in[177] ),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_1 _1351_ (.A(\grid_clb_1__1_.Q_in[178] ),
    .Y(_0366_));
 sky130_fd_sc_hd__inv_1 _1352_ (.A(\grid_clb_1__1_.Q_in[179] ),
    .Y(_0367_));
 sky130_fd_sc_hd__inv_1 _1353_ (.A(\grid_clb_1__1_.Q_in[172] ),
    .Y(_0360_));
 sky130_fd_sc_hd__inv_1 _1354_ (.A(\grid_clb_1__1_.Q_in[173] ),
    .Y(_0361_));
 sky130_fd_sc_hd__inv_1 _1355_ (.A(\grid_clb_1__1_.Q_in[174] ),
    .Y(_0362_));
 sky130_fd_sc_hd__inv_1 _1356_ (.A(\grid_clb_1__1_.Q_in[175] ),
    .Y(_0363_));
 sky130_fd_sc_hd__inv_1 _1357_ (.A(\grid_clb_1__1_.Q_in[184] ),
    .Y(_0372_));
 sky130_fd_sc_hd__inv_1 _1358_ (.A(\grid_clb_1__1_.Q_in[185] ),
    .Y(_0373_));
 sky130_fd_sc_hd__inv_1 _1359_ (.A(\grid_clb_1__1_.Q_in[186] ),
    .Y(_0374_));
 sky130_fd_sc_hd__inv_1 _1360_ (.A(\grid_clb_1__1_.Q_in[187] ),
    .Y(_0375_));
 sky130_fd_sc_hd__inv_1 _1361_ (.A(\grid_clb_1__1_.Q_in[180] ),
    .Y(_0368_));
 sky130_fd_sc_hd__inv_1 _1362_ (.A(\grid_clb_1__1_.Q_in[181] ),
    .Y(_0369_));
 sky130_fd_sc_hd__inv_1 _1363_ (.A(\grid_clb_1__1_.Q_in[182] ),
    .Y(_0370_));
 sky130_fd_sc_hd__inv_1 _1364_ (.A(\grid_clb_1__1_.Q_in[183] ),
    .Y(_0371_));
 sky130_fd_sc_hd__inv_1 _1365_ (.A(\grid_clb_1__1_.Q_in[192] ),
    .Y(_0380_));
 sky130_fd_sc_hd__inv_1 _1366_ (.A(\grid_clb_1__1_.Q_in[193] ),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_1 _1367_ (.A(\grid_clb_1__1_.Q_in[194] ),
    .Y(_0382_));
 sky130_fd_sc_hd__inv_1 _1368_ (.A(\grid_clb_1__1_.Q_in[195] ),
    .Y(_0383_));
 sky130_fd_sc_hd__inv_1 _1369_ (.A(\grid_clb_1__1_.Q_in[188] ),
    .Y(_0376_));
 sky130_fd_sc_hd__inv_1 _1370_ (.A(\grid_clb_1__1_.Q_in[189] ),
    .Y(_0377_));
 sky130_fd_sc_hd__inv_1 _1371_ (.A(\grid_clb_1__1_.Q_in[190] ),
    .Y(_0378_));
 sky130_fd_sc_hd__inv_1 _1372_ (.A(\grid_clb_1__1_.Q_in[191] ),
    .Y(_0379_));
 sky130_fd_sc_hd__inv_1 _1373_ (.A(\grid_clb_1__1_.Q_in[200] ),
    .Y(_0388_));
 sky130_fd_sc_hd__inv_1 _1374_ (.A(\grid_clb_1__1_.Q_in[201] ),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_1 _1375_ (.A(\grid_clb_1__1_.Q_in[202] ),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_1 _1376_ (.A(\grid_clb_1__1_.Q_in[203] ),
    .Y(_0391_));
 sky130_fd_sc_hd__inv_1 _1377_ (.A(\grid_clb_1__1_.Q_in[196] ),
    .Y(_0384_));
 sky130_fd_sc_hd__inv_1 _1378_ (.A(\grid_clb_1__1_.Q_in[197] ),
    .Y(_0385_));
 sky130_fd_sc_hd__inv_1 _1379_ (.A(\grid_clb_1__1_.Q_in[198] ),
    .Y(_0386_));
 sky130_fd_sc_hd__inv_1 _1380_ (.A(\grid_clb_1__1_.Q_in[199] ),
    .Y(_0387_));
 sky130_fd_sc_hd__inv_1 _1381_ (.A(\sb_0__0_.Q_in[62] ),
    .Y(_0406_));
 sky130_fd_sc_hd__inv_1 _1382_ (.A(\sb_0__0_.Q_in[61] ),
    .Y(_0405_));
 sky130_fd_sc_hd__inv_1 _1383_ (.A(\sb_0__0_.Q_in[60] ),
    .Y(_0404_));
 sky130_fd_sc_hd__inv_1 _1384_ (.A(\sb_0__0_.Q_in[65] ),
    .Y(_0409_));
 sky130_fd_sc_hd__inv_1 _1385_ (.A(\sb_0__0_.Q_in[64] ),
    .Y(_0408_));
 sky130_fd_sc_hd__inv_1 _1386_ (.A(\sb_0__0_.Q_in[63] ),
    .Y(_0407_));
 sky130_fd_sc_hd__inv_1 _1387_ (.A(\sb_0__0_.Q_in[56] ),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_1 _1388_ (.A(\sb_0__0_.Q_in[55] ),
    .Y(_0399_));
 sky130_fd_sc_hd__inv_1 _1389_ (.A(\sb_0__0_.Q_in[54] ),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_1 _1390_ (.A(\sb_0__0_.Q_in[59] ),
    .Y(_0403_));
 sky130_fd_sc_hd__inv_1 _1391_ (.A(\sb_0__0_.Q_in[58] ),
    .Y(_0402_));
 sky130_fd_sc_hd__inv_1 _1392_ (.A(\sb_0__0_.Q_in[57] ),
    .Y(_0401_));
 sky130_fd_sc_hd__inv_1 _1393_ (.A(\sb_0__0_.Q_in[42] ),
    .Y(_0412_));
 sky130_fd_sc_hd__inv_1 _1394_ (.A(\sb_0__0_.Q_in[41] ),
    .Y(_0411_));
 sky130_fd_sc_hd__inv_1 _1395_ (.A(\sb_0__0_.Q_in[40] ),
    .Y(_0410_));
 sky130_fd_sc_hd__inv_1 _1396_ (.A(\sb_0__0_.Q_in[45] ),
    .Y(_0415_));
 sky130_fd_sc_hd__inv_1 _1397_ (.A(\sb_0__0_.Q_in[44] ),
    .Y(_0414_));
 sky130_fd_sc_hd__inv_1 _1398_ (.A(\sb_0__0_.Q_in[43] ),
    .Y(_0413_));
 sky130_fd_sc_hd__inv_1 _1399_ (.A(\sb_0__0_.Q_in[36] ),
    .Y(_0394_));
 sky130_fd_sc_hd__inv_1 _1400_ (.A(\sb_0__0_.Q_in[35] ),
    .Y(_0393_));
 sky130_fd_sc_hd__inv_1 _1401_ (.A(\sb_0__0_.Q_in[34] ),
    .Y(_0392_));
 sky130_fd_sc_hd__inv_1 _1402_ (.A(\sb_0__0_.Q_in[39] ),
    .Y(_0397_));
 sky130_fd_sc_hd__inv_1 _1403_ (.A(\sb_0__0_.Q_in[38] ),
    .Y(_0396_));
 sky130_fd_sc_hd__inv_1 _1404_ (.A(\sb_0__0_.Q_in[37] ),
    .Y(_0395_));
 sky130_fd_sc_hd__inv_1 _1405_ (.A(\sb_0__0_.Q_in[18] ),
    .Y(_0424_));
 sky130_fd_sc_hd__inv_1 _1406_ (.A(\sb_0__0_.Q_in[17] ),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_1 _1407_ (.A(\sb_0__0_.Q_in[16] ),
    .Y(_0422_));
 sky130_fd_sc_hd__inv_1 _1408_ (.A(\sb_0__0_.Q_in[21] ),
    .Y(_0427_));
 sky130_fd_sc_hd__inv_1 _1409_ (.A(\sb_0__0_.Q_in[20] ),
    .Y(_0426_));
 sky130_fd_sc_hd__inv_1 _1410_ (.A(\sb_0__0_.Q_in[19] ),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_1 _1411_ (.A(\sb_0__0_.Q_in[2] ),
    .Y(_0418_));
 sky130_fd_sc_hd__inv_1 _1412_ (.A(\sb_0__0_.Q_in[1] ),
    .Y(_0417_));
 sky130_fd_sc_hd__inv_1 _1413_ (.A(\sb_0__0_.Q_in[0] ),
    .Y(_0416_));
 sky130_fd_sc_hd__inv_1 _1414_ (.A(\sb_0__0_.Q_in[5] ),
    .Y(_0421_));
 sky130_fd_sc_hd__inv_1 _1415_ (.A(\sb_0__0_.Q_in[4] ),
    .Y(_0420_));
 sky130_fd_sc_hd__inv_1 _1416_ (.A(\sb_0__0_.Q_in[3] ),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_1 _1417_ (.A(\sb_0__1_.Q_in[58] ),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_1 _1418_ (.A(\sb_0__1_.Q_in[57] ),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_1 _1419_ (.A(\sb_0__1_.Q_in[56] ),
    .Y(_0434_));
 sky130_fd_sc_hd__inv_1 _1420_ (.A(\sb_0__1_.Q_in[61] ),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_1 _1421_ (.A(\sb_0__1_.Q_in[60] ),
    .Y(_0438_));
 sky130_fd_sc_hd__inv_1 _1422_ (.A(\sb_0__1_.Q_in[59] ),
    .Y(_0437_));
 sky130_fd_sc_hd__inv_1 _1423_ (.A(\sb_0__1_.Q_in[42] ),
    .Y(_0442_));
 sky130_fd_sc_hd__inv_1 _1424_ (.A(\sb_0__1_.Q_in[41] ),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_1 _1425_ (.A(\sb_0__1_.Q_in[40] ),
    .Y(_0440_));
 sky130_fd_sc_hd__inv_1 _1426_ (.A(\sb_0__1_.Q_in[45] ),
    .Y(_0445_));
 sky130_fd_sc_hd__inv_1 _1427_ (.A(\sb_0__1_.Q_in[44] ),
    .Y(_0444_));
 sky130_fd_sc_hd__inv_1 _1428_ (.A(\sb_0__1_.Q_in[43] ),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_1 _1429_ (.A(\sb_0__1_.Q_in[36] ),
    .Y(_0430_));
 sky130_fd_sc_hd__inv_1 _1430_ (.A(\sb_0__1_.Q_in[35] ),
    .Y(_0429_));
 sky130_fd_sc_hd__inv_1 _1431_ (.A(\sb_0__1_.Q_in[34] ),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_1 _1432_ (.A(\sb_0__1_.Q_in[39] ),
    .Y(_0433_));
 sky130_fd_sc_hd__inv_1 _1433_ (.A(\sb_0__1_.Q_in[38] ),
    .Y(_0432_));
 sky130_fd_sc_hd__inv_1 _1434_ (.A(\sb_0__1_.Q_in[37] ),
    .Y(_0431_));
 sky130_fd_sc_hd__inv_1 _1435_ (.A(\sb_0__1_.Q_in[18] ),
    .Y(_0448_));
 sky130_fd_sc_hd__inv_1 _1436_ (.A(\sb_0__1_.Q_in[17] ),
    .Y(_0447_));
 sky130_fd_sc_hd__inv_1 _1437_ (.A(\sb_0__1_.Q_in[16] ),
    .Y(_0446_));
 sky130_fd_sc_hd__inv_1 _1438_ (.A(\sb_0__1_.Q_in[21] ),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_1 _1439_ (.A(\sb_0__1_.Q_in[20] ),
    .Y(_0450_));
 sky130_fd_sc_hd__inv_1 _1440_ (.A(\sb_0__1_.Q_in[19] ),
    .Y(_0449_));
 sky130_fd_sc_hd__inv_1 _1441_ (.A(\sb_1__0_.Q_in[66] ),
    .Y(_0466_));
 sky130_fd_sc_hd__inv_1 _1442_ (.A(\sb_1__0_.Q_in[65] ),
    .Y(_0465_));
 sky130_fd_sc_hd__inv_1 _1443_ (.A(\sb_1__0_.Q_in[64] ),
    .Y(_0464_));
 sky130_fd_sc_hd__inv_1 _1444_ (.A(\sb_1__0_.Q_in[69] ),
    .Y(_0469_));
 sky130_fd_sc_hd__inv_1 _1445_ (.A(\sb_1__0_.Q_in[68] ),
    .Y(_0468_));
 sky130_fd_sc_hd__inv_1 _1446_ (.A(\sb_1__0_.Q_in[67] ),
    .Y(_0467_));
 sky130_fd_sc_hd__inv_1 _1447_ (.A(\sb_1__0_.Q_in[60] ),
    .Y(_0460_));
 sky130_fd_sc_hd__inv_1 _1448_ (.A(\sb_1__0_.Q_in[59] ),
    .Y(_0459_));
 sky130_fd_sc_hd__inv_1 _1449_ (.A(\sb_1__0_.Q_in[58] ),
    .Y(_0458_));
 sky130_fd_sc_hd__inv_1 _1450_ (.A(\sb_1__0_.Q_in[63] ),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_1 _1451_ (.A(\sb_1__0_.Q_in[62] ),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_1 _1452_ (.A(\sb_1__0_.Q_in[61] ),
    .Y(_0461_));
 sky130_fd_sc_hd__inv_1 _1453_ (.A(\sb_1__0_.Q_in[46] ),
    .Y(_0472_));
 sky130_fd_sc_hd__inv_1 _1454_ (.A(\sb_1__0_.Q_in[45] ),
    .Y(_0471_));
 sky130_fd_sc_hd__inv_1 _1455_ (.A(\sb_1__0_.Q_in[44] ),
    .Y(_0470_));
 sky130_fd_sc_hd__inv_1 _1456_ (.A(\sb_1__0_.Q_in[49] ),
    .Y(_0475_));
 sky130_fd_sc_hd__inv_1 _1457_ (.A(\sb_1__0_.Q_in[48] ),
    .Y(_0474_));
 sky130_fd_sc_hd__inv_1 _1458_ (.A(\sb_1__0_.Q_in[47] ),
    .Y(_0473_));
 sky130_fd_sc_hd__inv_1 _1459_ (.A(\sb_1__0_.Q_in[40] ),
    .Y(_0454_));
 sky130_fd_sc_hd__inv_1 _1460_ (.A(\sb_1__0_.Q_in[39] ),
    .Y(_0453_));
 sky130_fd_sc_hd__inv_1 _1461_ (.A(\sb_1__0_.Q_in[38] ),
    .Y(_0452_));
 sky130_fd_sc_hd__inv_1 _1462_ (.A(\sb_1__0_.Q_in[43] ),
    .Y(_0457_));
 sky130_fd_sc_hd__inv_1 _1463_ (.A(\sb_1__0_.Q_in[42] ),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_1 _1464_ (.A(\sb_1__0_.Q_in[41] ),
    .Y(_0455_));
 sky130_fd_sc_hd__inv_1 _1465_ (.A(\sb_1__0_.Q_in[24] ),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_1 _1466_ (.A(\sb_1__0_.Q_in[23] ),
    .Y(_0483_));
 sky130_fd_sc_hd__inv_1 _1467_ (.A(\sb_1__0_.Q_in[22] ),
    .Y(_0482_));
 sky130_fd_sc_hd__inv_1 _1468_ (.A(\sb_1__0_.Q_in[27] ),
    .Y(_0487_));
 sky130_fd_sc_hd__inv_1 _1469_ (.A(\sb_1__0_.Q_in[26] ),
    .Y(_0486_));
 sky130_fd_sc_hd__inv_1 _1470_ (.A(\sb_1__0_.Q_in[25] ),
    .Y(_0485_));
 sky130_fd_sc_hd__inv_1 _1471_ (.A(\sb_1__0_.Q_in[8] ),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_1 _1472_ (.A(\sb_1__0_.Q_in[7] ),
    .Y(_0489_));
 sky130_fd_sc_hd__inv_1 _1473_ (.A(\sb_1__0_.Q_in[6] ),
    .Y(_0488_));
 sky130_fd_sc_hd__inv_1 _1474_ (.A(\sb_1__0_.Q_in[11] ),
    .Y(_0493_));
 sky130_fd_sc_hd__inv_1 _1475_ (.A(\sb_1__0_.Q_in[10] ),
    .Y(_0492_));
 sky130_fd_sc_hd__inv_1 _1476_ (.A(\sb_1__0_.Q_in[9] ),
    .Y(_0491_));
 sky130_fd_sc_hd__inv_1 _1477_ (.A(\sb_1__0_.Q_in[2] ),
    .Y(_0478_));
 sky130_fd_sc_hd__inv_1 _1478_ (.A(\sb_1__0_.Q_in[1] ),
    .Y(_0477_));
 sky130_fd_sc_hd__inv_1 _1479_ (.A(\sb_1__0_.Q_in[0] ),
    .Y(_0476_));
 sky130_fd_sc_hd__inv_1 _1480_ (.A(\sb_1__0_.Q_in[5] ),
    .Y(_0481_));
 sky130_fd_sc_hd__inv_1 _1481_ (.A(\sb_1__0_.Q_in[4] ),
    .Y(_0480_));
 sky130_fd_sc_hd__inv_1 _1482_ (.A(\sb_1__0_.Q_in[3] ),
    .Y(_0479_));
 sky130_fd_sc_hd__inv_1 _1483_ (.A(\sb_1__1_.Q_in[52] ),
    .Y(_0514_));
 sky130_fd_sc_hd__inv_1 _1484_ (.A(\sb_1__1_.Q_in[51] ),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_1 _1485_ (.A(\sb_1__1_.Q_in[50] ),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_1 _1486_ (.A(\sb_1__1_.Q_in[55] ),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_1 _1487_ (.A(\sb_1__1_.Q_in[54] ),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_1 _1488_ (.A(\sb_1__1_.Q_in[53] ),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_1 _1489_ (.A(\sb_1__1_.Q_in[36] ),
    .Y(_0508_));
 sky130_fd_sc_hd__inv_1 _1490_ (.A(\sb_1__1_.Q_in[35] ),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_1 _1491_ (.A(\sb_1__1_.Q_in[34] ),
    .Y(_0506_));
 sky130_fd_sc_hd__inv_1 _1492_ (.A(\sb_1__1_.Q_in[39] ),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_1 _1493_ (.A(\sb_1__1_.Q_in[38] ),
    .Y(_0510_));
 sky130_fd_sc_hd__inv_1 _1494_ (.A(\sb_1__1_.Q_in[37] ),
    .Y(_0509_));
 sky130_fd_sc_hd__inv_1 _1495_ (.A(\sb_1__1_.Q_in[18] ),
    .Y(_0502_));
 sky130_fd_sc_hd__inv_1 _1496_ (.A(\sb_1__1_.Q_in[17] ),
    .Y(_0501_));
 sky130_fd_sc_hd__inv_1 _1497_ (.A(\sb_1__1_.Q_in[16] ),
    .Y(_0500_));
 sky130_fd_sc_hd__inv_1 _1498_ (.A(\sb_1__1_.Q_in[21] ),
    .Y(_0505_));
 sky130_fd_sc_hd__inv_1 _1499_ (.A(\sb_1__1_.Q_in[20] ),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_1 _1500_ (.A(\sb_1__1_.Q_in[19] ),
    .Y(_0503_));
 sky130_fd_sc_hd__inv_1 _1501_ (.A(\sb_1__1_.Q_in[2] ),
    .Y(_0496_));
 sky130_fd_sc_hd__inv_1 _1502_ (.A(\sb_1__1_.Q_in[1] ),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_1 _1503_ (.A(\sb_1__1_.Q_in[0] ),
    .Y(_0494_));
 sky130_fd_sc_hd__inv_1 _1504_ (.A(\sb_1__1_.Q_in[5] ),
    .Y(_0499_));
 sky130_fd_sc_hd__inv_1 _1505_ (.A(\sb_1__1_.Q_in[4] ),
    .Y(_0498_));
 sky130_fd_sc_hd__inv_1 _1506_ (.A(\sb_1__1_.Q_in[3] ),
    .Y(_0497_));
 sky130_fd_sc_hd__inv_1 _1507_ (.A(\cbx_1__0_.Q_in[62] ),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_1 _1508_ (.A(\cbx_1__0_.Q_in[61] ),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_1 _1509_ (.A(\cbx_1__0_.Q_in[60] ),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_1 _1510_ (.A(\cbx_1__0_.Q_in[65] ),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_1 _1511_ (.A(\cbx_1__0_.Q_in[64] ),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_1 _1512_ (.A(\cbx_1__0_.Q_in[63] ),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_1 _1513_ (.A(\cbx_1__0_.Q_in[56] ),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_1 _1514_ (.A(\cbx_1__0_.Q_in[55] ),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_1 _1515_ (.A(\cbx_1__0_.Q_in[54] ),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_1 _1516_ (.A(\cbx_1__0_.Q_in[59] ),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_1 _1517_ (.A(\cbx_1__0_.Q_in[58] ),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_1 _1518_ (.A(\cbx_1__0_.Q_in[57] ),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_1 _1519_ (.A(\cbx_1__0_.Q_in[50] ),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_1 _1520_ (.A(\cbx_1__0_.Q_in[49] ),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_1 _1521_ (.A(\cbx_1__0_.Q_in[48] ),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_1 _1522_ (.A(\cbx_1__0_.Q_in[53] ),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_1 _1523_ (.A(\cbx_1__0_.Q_in[52] ),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_1 _1524_ (.A(\cbx_1__0_.Q_in[51] ),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_1 _1525_ (.A(\cbx_1__0_.Q_in[44] ),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_1 _1526_ (.A(\cbx_1__0_.Q_in[43] ),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_1 _1527_ (.A(\cbx_1__0_.Q_in[42] ),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_1 _1528_ (.A(\cbx_1__0_.Q_in[47] ),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_1 _1529_ (.A(\cbx_1__0_.Q_in[46] ),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_1 _1530_ (.A(\cbx_1__0_.Q_in[45] ),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_1 _1531_ (.A(\cbx_1__0_.Q_in[38] ),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_1 _1532_ (.A(\cbx_1__0_.Q_in[37] ),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_1 _1533_ (.A(\cbx_1__0_.Q_in[36] ),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_1 _1534_ (.A(\cbx_1__0_.Q_in[41] ),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_1 _1535_ (.A(\cbx_1__0_.Q_in[40] ),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_1 _1536_ (.A(\cbx_1__0_.Q_in[39] ),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_1 _1537_ (.A(\cbx_1__0_.Q_in[32] ),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_1 _1538_ (.A(\cbx_1__0_.Q_in[31] ),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_1 _1539_ (.A(\cbx_1__0_.Q_in[30] ),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_1 _1540_ (.A(\cbx_1__0_.Q_in[35] ),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_1 _1541_ (.A(\cbx_1__0_.Q_in[34] ),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_1 _1542_ (.A(\cbx_1__0_.Q_in[33] ),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_1 _1543_ (.A(\cbx_1__0_.Q_in[26] ),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_1 _1544_ (.A(\cbx_1__0_.Q_in[25] ),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_1 _1545_ (.A(\cbx_1__0_.Q_in[24] ),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_1 _1546_ (.A(\cbx_1__0_.Q_in[29] ),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_1 _1547_ (.A(\cbx_1__0_.Q_in[28] ),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_1 _1548_ (.A(\cbx_1__0_.Q_in[27] ),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_1 _1549_ (.A(\cbx_1__0_.Q_in[20] ),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_1 _1550_ (.A(\cbx_1__0_.Q_in[19] ),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_1 _1551_ (.A(\cbx_1__0_.Q_in[18] ),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_1 _1552_ (.A(\cbx_1__0_.Q_in[23] ),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_1 _1553_ (.A(\cbx_1__0_.Q_in[22] ),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_1 _1554_ (.A(\cbx_1__0_.Q_in[21] ),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_1 _1555_ (.A(\cbx_1__0_.Q_in[8] ),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_1 _1556_ (.A(\cbx_1__0_.Q_in[7] ),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_1 _1557_ (.A(\cbx_1__0_.Q_in[6] ),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_1 _1558_ (.A(\cbx_1__0_.Q_in[11] ),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_1 _1559_ (.A(\cbx_1__0_.Q_in[10] ),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_1 _1560_ (.A(\cbx_1__0_.Q_in[9] ),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_1 _1561_ (.A(\cbx_1__0_.Q_in[2] ),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_1 _1562_ (.A(\cbx_1__0_.Q_in[1] ),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_1 _1563_ (.A(\cbx_1__0_.Q_in[0] ),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_1 _1564_ (.A(\cbx_1__0_.Q_in[5] ),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_1 _1565_ (.A(\cbx_1__0_.Q_in[4] ),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_1 _1566_ (.A(\cbx_1__0_.Q_in[3] ),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_1 _1567_ (.A(\cbx_1__1_.Q_in[62] ),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_1 _1568_ (.A(\cbx_1__1_.Q_in[61] ),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_1 _1569_ (.A(\cbx_1__1_.Q_in[60] ),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_1 _1570_ (.A(\cbx_1__1_.Q_in[65] ),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_1 _1571_ (.A(\cbx_1__1_.Q_in[64] ),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_1 _1572_ (.A(\cbx_1__1_.Q_in[63] ),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_1 _1573_ (.A(\cbx_1__1_.Q_in[56] ),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_1 _1574_ (.A(\cbx_1__1_.Q_in[55] ),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_1 _1575_ (.A(\cbx_1__1_.Q_in[54] ),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_1 _1576_ (.A(\cbx_1__1_.Q_in[59] ),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_1 _1577_ (.A(\cbx_1__1_.Q_in[58] ),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_1 _1578_ (.A(\cbx_1__1_.Q_in[57] ),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_1 _1579_ (.A(\cbx_1__1_.Q_in[50] ),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_1 _1580_ (.A(\cbx_1__1_.Q_in[49] ),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_1 _1581_ (.A(\cbx_1__1_.Q_in[48] ),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_1 _1582_ (.A(\cbx_1__1_.Q_in[53] ),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_1 _1583_ (.A(\cbx_1__1_.Q_in[52] ),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_1 _1584_ (.A(\cbx_1__1_.Q_in[51] ),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_1 _1585_ (.A(\cbx_1__1_.Q_in[44] ),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_1 _1586_ (.A(\cbx_1__1_.Q_in[43] ),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_1 _1587_ (.A(\cbx_1__1_.Q_in[42] ),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_1 _1588_ (.A(\cbx_1__1_.Q_in[47] ),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_1 _1589_ (.A(\cbx_1__1_.Q_in[46] ),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_1 _1590_ (.A(\cbx_1__1_.Q_in[45] ),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_1 _1591_ (.A(\cbx_1__1_.Q_in[38] ),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_1 _1592_ (.A(\cbx_1__1_.Q_in[37] ),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_1 _1593_ (.A(\cbx_1__1_.Q_in[36] ),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_1 _1594_ (.A(\cbx_1__1_.Q_in[41] ),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_1 _1595_ (.A(\cbx_1__1_.Q_in[40] ),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_1 _1596_ (.A(\cbx_1__1_.Q_in[39] ),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_1 _1597_ (.A(\cbx_1__1_.Q_in[32] ),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_1 _1598_ (.A(\cbx_1__1_.Q_in[31] ),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_1 _1599_ (.A(\cbx_1__1_.Q_in[30] ),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_1 _1600_ (.A(\cbx_1__1_.Q_in[35] ),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_1 _1601_ (.A(\cbx_1__1_.Q_in[34] ),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_1 _1602_ (.A(\cbx_1__1_.Q_in[33] ),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_1 _1603_ (.A(\cbx_1__1_.Q_in[26] ),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_1 _1604_ (.A(\cbx_1__1_.Q_in[25] ),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_1 _1605_ (.A(\cbx_1__1_.Q_in[24] ),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_1 _1606_ (.A(\cbx_1__1_.Q_in[29] ),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_1 _1607_ (.A(\cbx_1__1_.Q_in[28] ),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_1 _1608_ (.A(\cbx_1__1_.Q_in[27] ),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_1 _1609_ (.A(\cbx_1__1_.Q_in[20] ),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_1 _1610_ (.A(\cbx_1__1_.Q_in[19] ),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_1 _1611_ (.A(\cbx_1__1_.Q_in[18] ),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_1 _1612_ (.A(\cbx_1__1_.Q_in[23] ),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_1 _1613_ (.A(\cbx_1__1_.Q_in[22] ),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_1 _1614_ (.A(\cbx_1__1_.Q_in[21] ),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_1 _1615_ (.A(\cbx_1__1_.Q_in[14] ),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_1 _1616_ (.A(\cbx_1__1_.Q_in[13] ),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_1 _1617_ (.A(\cbx_1__1_.Q_in[12] ),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_1 _1618_ (.A(\cbx_1__1_.Q_in[17] ),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_1 _1619_ (.A(\cbx_1__1_.Q_in[16] ),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_1 _1620_ (.A(\cbx_1__1_.Q_in[15] ),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_1 _1621_ (.A(\cbx_1__1_.Q_in[8] ),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_1 _1622_ (.A(\cbx_1__1_.Q_in[7] ),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_1 _1623_ (.A(\cbx_1__1_.Q_in[6] ),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_1 _1624_ (.A(\cbx_1__1_.Q_in[11] ),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_1 _1625_ (.A(\cbx_1__1_.Q_in[10] ),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_1 _1626_ (.A(\cbx_1__1_.Q_in[9] ),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_1 _1627_ (.A(\cbx_1__1_.Q_in[2] ),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_1 _1628_ (.A(\cbx_1__1_.Q_in[1] ),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_1 _1629_ (.A(\cbx_1__1_.Q_in[0] ),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_1 _1630_ (.A(\cbx_1__1_.Q_in[5] ),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_1 _1631_ (.A(\cbx_1__1_.Q_in[4] ),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_1 _1632_ (.A(\cbx_1__1_.Q_in[3] ),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_1 _1633_ (.A(\cby_0__1_.Q_in[56] ),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_1 _1634_ (.A(\cby_0__1_.Q_in[55] ),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_1 _1635_ (.A(\cby_0__1_.Q_in[54] ),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_1 _1636_ (.A(\cby_0__1_.Q_in[59] ),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_1 _1637_ (.A(\cby_0__1_.Q_in[58] ),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_1 _1638_ (.A(\cby_0__1_.Q_in[57] ),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_1 _1639_ (.A(\cby_0__1_.Q_in[50] ),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_1 _1640_ (.A(\cby_0__1_.Q_in[49] ),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_1 _1641_ (.A(\cby_0__1_.Q_in[48] ),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_1 _1642_ (.A(\cby_0__1_.Q_in[53] ),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_1 _1643_ (.A(\cby_0__1_.Q_in[52] ),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_1 _1644_ (.A(\cby_0__1_.Q_in[51] ),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_1 _1645_ (.A(\cby_0__1_.Q_in[44] ),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_1 _1646_ (.A(\cby_0__1_.Q_in[43] ),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_1 _1647_ (.A(\cby_0__1_.Q_in[42] ),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_1 _1648_ (.A(\cby_0__1_.Q_in[47] ),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_1 _1649_ (.A(\cby_0__1_.Q_in[46] ),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_1 _1650_ (.A(\cby_0__1_.Q_in[45] ),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_1 _1651_ (.A(\cby_0__1_.Q_in[38] ),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_1 _1652_ (.A(\cby_0__1_.Q_in[37] ),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_1 _1653_ (.A(\cby_0__1_.Q_in[36] ),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_1 _1654_ (.A(\cby_0__1_.Q_in[41] ),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_1 _1655_ (.A(\cby_0__1_.Q_in[40] ),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_1 _1656_ (.A(\cby_0__1_.Q_in[39] ),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_1 _1657_ (.A(\cby_0__1_.Q_in[32] ),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_1 _1658_ (.A(\cby_0__1_.Q_in[31] ),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_1 _1659_ (.A(\cby_0__1_.Q_in[30] ),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_1 _1660_ (.A(\cby_0__1_.Q_in[35] ),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_1 _1661_ (.A(\cby_0__1_.Q_in[34] ),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_1 _1662_ (.A(\cby_0__1_.Q_in[33] ),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_1 _1663_ (.A(\cby_0__1_.Q_in[26] ),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_1 _1664_ (.A(\cby_0__1_.Q_in[25] ),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_1 _1665_ (.A(\cby_0__1_.Q_in[24] ),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_1 _1666_ (.A(\cby_0__1_.Q_in[29] ),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_1 _1667_ (.A(\cby_0__1_.Q_in[28] ),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_1 _1668_ (.A(\cby_0__1_.Q_in[27] ),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_1 _1669_ (.A(\cby_0__1_.Q_in[20] ),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_1 _1670_ (.A(\cby_0__1_.Q_in[19] ),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_1 _1671_ (.A(\cby_0__1_.Q_in[18] ),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_1 _1672_ (.A(\cby_0__1_.Q_in[23] ),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_1 _1673_ (.A(\cby_0__1_.Q_in[22] ),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_1 _1674_ (.A(\cby_0__1_.Q_in[21] ),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_1 _1675_ (.A(\cby_0__1_.Q_in[14] ),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_1 _1676_ (.A(\cby_0__1_.Q_in[13] ),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_1 _1677_ (.A(\cby_0__1_.Q_in[12] ),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_1 _1678_ (.A(\cby_0__1_.Q_in[17] ),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_1 _1679_ (.A(\cby_0__1_.Q_in[16] ),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_1 _1680_ (.A(\cby_0__1_.Q_in[15] ),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_1 _1681_ (.A(\cby_0__1_.Q_in[8] ),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_1 _1682_ (.A(\cby_0__1_.Q_in[7] ),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_1 _1683_ (.A(\cby_0__1_.Q_in[6] ),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_1 _1684_ (.A(\cby_0__1_.Q_in[11] ),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_1 _1685_ (.A(\cby_0__1_.Q_in[10] ),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_1 _1686_ (.A(\cby_0__1_.Q_in[9] ),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_1 _1687_ (.A(\cby_0__1_.Q_in[2] ),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_1 _1688_ (.A(\cby_0__1_.Q_in[1] ),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_1 _1689_ (.A(\cby_0__1_.Q_in[0] ),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_1 _1690_ (.A(\cby_0__1_.Q_in[5] ),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_1 _1691_ (.A(\cby_0__1_.Q_in[4] ),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_1 _1692_ (.A(\cby_0__1_.Q_in[3] ),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_1 _1693_ (.A(\cby_1__1_.Q_in[62] ),
    .Y(_0248_));
 sky130_fd_sc_hd__inv_1 _1694_ (.A(\cby_1__1_.Q_in[61] ),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_1 _1695_ (.A(\cby_1__1_.Q_in[60] ),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_1 _1696_ (.A(\cby_1__1_.Q_in[65] ),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_1 _1697_ (.A(\cby_1__1_.Q_in[64] ),
    .Y(_0250_));
 sky130_fd_sc_hd__inv_1 _1698_ (.A(\cby_1__1_.Q_in[63] ),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_1 _1699_ (.A(\cby_1__1_.Q_in[56] ),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_1 _1700_ (.A(\cby_1__1_.Q_in[55] ),
    .Y(_0241_));
 sky130_fd_sc_hd__inv_1 _1701_ (.A(\cby_1__1_.Q_in[54] ),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_1 _1702_ (.A(\cby_1__1_.Q_in[59] ),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_1 _1703_ (.A(\cby_1__1_.Q_in[58] ),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_1 _1704_ (.A(\cby_1__1_.Q_in[57] ),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_1 _1705_ (.A(\cby_1__1_.Q_in[50] ),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_1 _1706_ (.A(\cby_1__1_.Q_in[49] ),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_1 _1707_ (.A(\cby_1__1_.Q_in[48] ),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_1 _1708_ (.A(\cby_1__1_.Q_in[53] ),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_1 _1709_ (.A(\cby_1__1_.Q_in[52] ),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_1 _1710_ (.A(\cby_1__1_.Q_in[51] ),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_1 _1711_ (.A(\cby_1__1_.Q_in[44] ),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_1 _1712_ (.A(\cby_1__1_.Q_in[43] ),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_1 _1713_ (.A(\cby_1__1_.Q_in[42] ),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_1 _1714_ (.A(\cby_1__1_.Q_in[47] ),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_1 _1715_ (.A(\cby_1__1_.Q_in[46] ),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_1 _1716_ (.A(\cby_1__1_.Q_in[45] ),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_1 _1717_ (.A(\cby_1__1_.Q_in[38] ),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_1 _1718_ (.A(\cby_1__1_.Q_in[37] ),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_1 _1719_ (.A(\cby_1__1_.Q_in[36] ),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_1 _1720_ (.A(\cby_1__1_.Q_in[41] ),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_1 _1721_ (.A(\cby_1__1_.Q_in[40] ),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_1 _1722_ (.A(\cby_1__1_.Q_in[39] ),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_1 _1723_ (.A(\cby_1__1_.Q_in[32] ),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_1 _1724_ (.A(\cby_1__1_.Q_in[31] ),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_1 _1725_ (.A(\cby_1__1_.Q_in[30] ),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_1 _1726_ (.A(\cby_1__1_.Q_in[35] ),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_1 _1727_ (.A(\cby_1__1_.Q_in[34] ),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_1 _1728_ (.A(\cby_1__1_.Q_in[33] ),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_1 _1729_ (.A(\cby_1__1_.Q_in[26] ),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_1 _1730_ (.A(\cby_1__1_.Q_in[25] ),
    .Y(_0211_));
 sky130_fd_sc_hd__inv_1 _1731_ (.A(\cby_1__1_.Q_in[24] ),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_1 _1732_ (.A(\cby_1__1_.Q_in[29] ),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_1 _1733_ (.A(\cby_1__1_.Q_in[28] ),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_1 _1734_ (.A(\cby_1__1_.Q_in[27] ),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_1 _1735_ (.A(\cby_1__1_.Q_in[20] ),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_1 _1736_ (.A(\cby_1__1_.Q_in[19] ),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_1 _1737_ (.A(\cby_1__1_.Q_in[18] ),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_1 _1738_ (.A(\cby_1__1_.Q_in[23] ),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_1 _1739_ (.A(\cby_1__1_.Q_in[22] ),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_1 _1740_ (.A(\cby_1__1_.Q_in[21] ),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_1 _1741_ (.A(\cby_1__1_.Q_in[14] ),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_1 _1742_ (.A(\cby_1__1_.Q_in[13] ),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_1 _1743_ (.A(\cby_1__1_.Q_in[12] ),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_1 _1744_ (.A(\cby_1__1_.Q_in[17] ),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_1 _1745_ (.A(\cby_1__1_.Q_in[16] ),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_1 _1746_ (.A(\cby_1__1_.Q_in[15] ),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_1 _1747_ (.A(\cby_1__1_.Q_in[8] ),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_1 _1748_ (.A(\cby_1__1_.Q_in[7] ),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_1 _1749_ (.A(\cby_1__1_.Q_in[6] ),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_1 _1750_ (.A(\cby_1__1_.Q_in[11] ),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_1 _1751_ (.A(\cby_1__1_.Q_in[10] ),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_1 _1752_ (.A(\cby_1__1_.Q_in[9] ),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_1 _1753_ (.A(\cby_1__1_.Q_in[2] ),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_1 _1754_ (.A(\cby_1__1_.Q_in[1] ),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_1 _1755_ (.A(\cby_1__1_.Q_in[0] ),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_1 _1756_ (.A(\cby_1__1_.Q_in[5] ),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_1 _1757_ (.A(\cby_1__1_.Q_in[4] ),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_1 _1758_ (.A(\cby_1__1_.Q_in[3] ),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_1 _1759_ (.A(\grid_clb_1__1_.Q_in[75] ),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_1 _1760_ (.A(\grid_clb_1__1_.Q_in[17] ),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_1 _1761_ (.A(\grid_clb_1__1_.Q_in[16] ),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_1 _1762_ (.A(\grid_clb_1__1_.Q_in[18] ),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_1 _1763_ (.A(\grid_clb_1__1_.Q_in[36] ),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_1 _1764_ (.A(\grid_clb_1__1_.Q_in[35] ),
    .Y(_0255_));
 sky130_fd_sc_hd__inv_1 _1765_ (.A(\grid_clb_1__1_.Q_in[37] ),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_1 _1766_ (.A(\grid_clb_1__1_.Q_in[55] ),
    .Y(_0259_));
 sky130_fd_sc_hd__inv_1 _1767_ (.A(\grid_clb_1__1_.Q_in[54] ),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_1 _1768_ (.A(\grid_clb_1__1_.Q_in[56] ),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_1 _1769_ (.A(\grid_clb_1__1_.Q_in[74] ),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_1 _1770_ (.A(\grid_clb_1__1_.Q_in[73] ),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_1 _1771_ (.A(\grid_clb_1__1_.Q_in[80] ),
    .Y(_0268_));
 sky130_fd_sc_hd__inv_1 _1772_ (.A(\grid_clb_1__1_.Q_in[81] ),
    .Y(_0269_));
 sky130_fd_sc_hd__inv_1 _1773_ (.A(\grid_clb_1__1_.Q_in[82] ),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_1 _1774_ (.A(\grid_clb_1__1_.Q_in[83] ),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_1 _1775_ (.A(\grid_clb_1__1_.Q_in[76] ),
    .Y(_0264_));
 sky130_fd_sc_hd__inv_1 _1776_ (.A(\grid_clb_1__1_.Q_in[77] ),
    .Y(_0265_));
 sky130_fd_sc_hd__inv_1 _1777_ (.A(\grid_clb_1__1_.Q_in[78] ),
    .Y(_0266_));
 sky130_fd_sc_hd__inv_1 _1778_ (.A(\grid_clb_1__1_.Q_in[79] ),
    .Y(_0267_));
 sky130_fd_sc_hd__inv_1 _1779_ (.A(\grid_clb_1__1_.Q_in[88] ),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_1 _1780_ (.A(\grid_clb_1__1_.Q_in[89] ),
    .Y(_0277_));
 sky130_fd_sc_hd__inv_1 _1781_ (.A(\grid_clb_1__1_.Q_in[90] ),
    .Y(_0278_));
 sky130_fd_sc_hd__inv_1 _1782_ (.A(\grid_clb_1__1_.Q_in[91] ),
    .Y(_0279_));
 sky130_fd_sc_hd__inv_1 _1783_ (.A(\grid_clb_1__1_.Q_in[84] ),
    .Y(_0272_));
 sky130_fd_sc_hd__inv_1 _1784_ (.A(\grid_clb_1__1_.Q_in[85] ),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_1 _1785_ (.A(\grid_clb_1__1_.Q_in[86] ),
    .Y(_0274_));
 sky130_fd_sc_hd__inv_1 _1786_ (.A(\grid_clb_1__1_.Q_in[87] ),
    .Y(_0275_));
 sky130_fd_sc_hd__inv_1 _1787_ (.A(\grid_clb_1__1_.Q_in[96] ),
    .Y(_0284_));
 sky130_fd_sc_hd__inv_1 _1788_ (.A(\grid_clb_1__1_.Q_in[97] ),
    .Y(_0285_));
 sky130_fd_sc_hd__inv_1 _1789_ (.A(\grid_clb_1__1_.Q_in[98] ),
    .Y(_0286_));
 sky130_fd_sc_hd__inv_1 _1790_ (.A(\grid_clb_1__1_.Q_in[99] ),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_1 _1791_ (.A(\grid_clb_1__1_.Q_in[92] ),
    .Y(_0280_));
 sky130_fd_sc_hd__inv_1 _1792_ (.A(\grid_clb_1__1_.Q_in[93] ),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_1 _1793_ (.A(\grid_clb_1__1_.Q_in[94] ),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_1 _1794_ (.A(\grid_clb_1__1_.Q_in[95] ),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_1 _1795_ (.A(reset),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _1796_ (.A(set),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__conb_1 _1797_ (.HI(_0725_));
 sky130_fd_sc_hd__dfbbp_1 _1798_ (.CLK(clk),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_ff_0.DFFSRQ_0_.D ),
    .RESET_B(_0518_),
    .SET_B(_0519_),
    .Q(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ),
    .Q_N(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__dfbbp_1 _1799_ (.CLK(clk),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_ff_0.DFFSRQ_0_.D ),
    .RESET_B(_0518_),
    .SET_B(_0519_),
    .Q(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ),
    .Q_N(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__dfbbp_1 _1800_ (.CLK(clk),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_ff_0.DFFSRQ_0_.D ),
    .RESET_B(_0518_),
    .SET_B(_0519_),
    .Q(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ),
    .Q_N(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__dfbbp_1 _1801_ (.CLK(clk),
    .D(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_ff_0.DFFSRQ_0_.D ),
    .RESET_B(_0518_),
    .SET_B(_0519_),
    .Q(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_ff_0.DFFSRQ_0_.Q ),
    .Q_N(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.INVTX1_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.out ),
    .TE_B(_0000_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.out ),
    .TE_B(_0001_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.out ),
    .TE_B(_0002_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.out ),
    .TE_B(_0000_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_0001_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_0002_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0003_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0004_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0005_),
    .Z(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.out ),
    .TE_B(_0006_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.out ),
    .TE_B(_0007_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.out ),
    .TE_B(_0008_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.out ),
    .TE_B(_0006_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.out ),
    .TE_B(_0007_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.out ),
    .TE_B(_0008_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0009_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0010_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0011_),
    .Z(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_0012_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_0013_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_0014_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_0012_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_4_.out ),
    .TE_B(_0013_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_5_.out ),
    .TE_B(_0014_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0015_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0016_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0017_),
    .Z(\cbx_1__0_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_0018_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_0019_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.INVTX1_2_.out ),
    .TE_B(_0020_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.INVTX1_3_.out ),
    .TE_B(_0018_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.INVTX1_4_.out ),
    .TE_B(_0019_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0020_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0021_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0022_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0023_),
    .Z(\cbx_1__0_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.INVTX1_2_.out ),
    .TE_B(_0024_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.INVTX1_3_.out ),
    .TE_B(_0025_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_2_.out ),
    .TE_B(_0026_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_3_.out ),
    .TE_B(_0024_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_4_.out ),
    .TE_B(_0025_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0026_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_0_.out ),
    .TE_B(_0027_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_2.mux_l1_in_1_.out ),
    .TE_B(_0028_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0029_),
    .Z(\cbx_1__0_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_2_.out ),
    .TE_B(_0030_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_2.INVTX1_3_.out ),
    .TE_B(_0031_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.out ),
    .TE_B(_0032_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.out ),
    .TE_B(_0030_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_0031_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_0032_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_0_.out ),
    .TE_B(_0033_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_3.mux_l1_in_1_.out ),
    .TE_B(_0034_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0035_),
    .Z(\cbx_1__0_.mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.out ),
    .TE_B(_0036_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.out ),
    .TE_B(_0037_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.out ),
    .TE_B(_0038_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.out ),
    .TE_B(_0036_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.out ),
    .TE_B(_0037_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.out ),
    .TE_B(_0038_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_0_.out ),
    .TE_B(_0039_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_4.mux_l1_in_1_.out ),
    .TE_B(_0040_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0041_),
    .Z(\cbx_1__0_.mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.out ),
    .TE_B(_0042_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.out ),
    .TE_B(_0043_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.out ),
    .TE_B(_0044_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.out ),
    .TE_B(_0042_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_0043_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_0044_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_0_.out ),
    .TE_B(_0045_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_5.mux_l1_in_1_.out ),
    .TE_B(_0046_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0047_),
    .Z(\cbx_1__0_.mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_2_.out ),
    .TE_B(_0048_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_0049_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_0050_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_0048_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_4_.out ),
    .TE_B(_0049_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_5_.out ),
    .TE_B(_0050_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_0_.out ),
    .TE_B(_0051_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_6.mux_l1_in_1_.out ),
    .TE_B(_0052_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0053_),
    .Z(\cbx_1__0_.mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_2_.out ),
    .TE_B(_0054_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_3_.out ),
    .TE_B(_0055_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_4_.out ),
    .TE_B(_0056_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_0.INVTX1_5_.out ),
    .TE_B(_0054_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_1.INVTX1_4_.out ),
    .TE_B(_0055_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0056_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_0_.out ),
    .TE_B(_0057_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_top_ipin_7.mux_l1_in_1_.out ),
    .TE_B(_0058_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0059_),
    .Z(\cbx_1__0_.mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.out ),
    .TE_B(_0060_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.out ),
    .TE_B(_0061_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.out ),
    .TE_B(_0062_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.out ),
    .TE_B(_0060_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_0061_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_0062_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0063_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0064_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0065_),
    .Z(\cbx_1__1_.mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.out ),
    .TE_B(_0066_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.out ),
    .TE_B(_0067_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0068_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_0066_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_0067_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_0068_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0069_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0070_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0071_),
    .Z(\cbx_1__1_.mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0072_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_0073_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0074_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_0072_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_0073_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_0074_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_0_.out ),
    .TE_B(_0075_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.mux_l1_in_1_.out ),
    .TE_B(_0076_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0077_),
    .Z(\cbx_1__1_.mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0078_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_0079_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0080_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_3_.out ),
    .TE_B(_0078_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_4_.out ),
    .TE_B(_0079_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_5_.out ),
    .TE_B(_0080_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_0_.out ),
    .TE_B(_0081_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.mux_l1_in_1_.out ),
    .TE_B(_0082_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0083_),
    .Z(\cbx_1__1_.mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0084_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_3_.out ),
    .TE_B(_0085_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0086_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_3_.out ),
    .TE_B(_0084_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_4_.out ),
    .TE_B(_0085_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_5_.out ),
    .TE_B(_0086_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_0_.out ),
    .TE_B(_0087_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.mux_l1_in_1_.out ),
    .TE_B(_0088_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0089_),
    .Z(\cbx_1__1_.mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0090_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_3_.out ),
    .TE_B(_0091_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_2_.out ),
    .TE_B(_0092_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_3_.out ),
    .TE_B(_0090_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_4_.out ),
    .TE_B(_0091_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_5_.out ),
    .TE_B(_0092_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_0_.out ),
    .TE_B(_0093_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.mux_l1_in_1_.out ),
    .TE_B(_0094_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0095_),
    .Z(\cbx_1__1_.mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_2_.out ),
    .TE_B(_0096_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_3_.out ),
    .TE_B(_0097_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.out ),
    .TE_B(_0098_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.out ),
    .TE_B(_0096_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_0097_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_0.INVTX1_5_.out ),
    .TE_B(_0098_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_0_.out ),
    .TE_B(_0099_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_6.mux_l1_in_1_.out ),
    .TE_B(_0100_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0101_),
    .Z(\cbx_1__1_.mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.out ),
    .TE_B(_0102_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.out ),
    .TE_B(_0103_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.out ),
    .TE_B(_0104_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.out ),
    .TE_B(_0102_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_0103_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_0104_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_0_.out ),
    .TE_B(_0105_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_7.mux_l1_in_1_.out ),
    .TE_B(_0106_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0107_),
    .Z(\cbx_1__1_.mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0108_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_3_.out ),
    .TE_B(_0109_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_0110_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_5_.out ),
    .TE_B(_0108_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_0109_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_0110_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0111_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0112_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0113_),
    .Z(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0114_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_3_.out ),
    .TE_B(_0115_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_4_.out ),
    .TE_B(_0116_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_2.INVTX1_5_.out ),
    .TE_B(_0114_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_4_.out ),
    .TE_B(_0115_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_5_.out ),
    .TE_B(_0116_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0117_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0118_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0119_),
    .Z(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0120_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_3_.out ),
    .TE_B(_0121_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_4_.out ),
    .TE_B(_0122_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_3.INVTX1_5_.out ),
    .TE_B(_0120_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_4_.out ),
    .TE_B(_0121_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_5_.out ),
    .TE_B(_0122_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_0_.out ),
    .TE_B(_0123_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l1_in_1_.out ),
    .TE_B(_0124_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0125_),
    .Z(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .TE_B(_0126_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0127_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.out ),
    .TE_B(_0128_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_3_.out ),
    .TE_B(_0126_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_4_.out ),
    .TE_B(_0127_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_0128_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0129_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0130_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0131_),
    .Z(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .TE_B(_0132_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0133_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .TE_B(_0134_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.out ),
    .TE_B(_0132_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .TE_B(_0133_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.out ),
    .TE_B(_0134_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0135_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0136_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0137_),
    .Z(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .TE_B(_0138_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.out ),
    .TE_B(_0139_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_2_.out ),
    .TE_B(_0140_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .TE_B(_0138_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_4_.out ),
    .TE_B(_0139_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_5_.out ),
    .TE_B(_0140_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0141_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0142_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0143_),
    .Z(\cby_0__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_2_.out ),
    .TE_B(_0144_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .TE_B(_0145_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.INVTX1_2_.out ),
    .TE_B(_0146_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.INVTX1_3_.out ),
    .TE_B(_0144_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0145_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.INVTX1_5_.out ),
    .TE_B(_0146_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0147_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0148_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0149_),
    .Z(\cby_0__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.INVTX1_2_.out ),
    .TE_B(_0150_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.INVTX1_3_.out ),
    .TE_B(_0151_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_2.INVTX1_2_.out ),
    .TE_B(_0152_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_2.INVTX1_3_.out ),
    .TE_B(_0150_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0151_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_2.INVTX1_5_.out ),
    .TE_B(_0152_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_2.mux_l1_in_0_.out ),
    .TE_B(_0153_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_2.mux_l1_in_1_.out ),
    .TE_B(_0154_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0155_),
    .Z(\cby_0__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_2.INVTX1_2_.out ),
    .TE_B(_0156_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_2.INVTX1_3_.out ),
    .TE_B(_0157_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_2_.out ),
    .TE_B(_0158_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_3_.out ),
    .TE_B(_0156_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_4_.out ),
    .TE_B(_0157_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_5_.out ),
    .TE_B(_0158_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.mux_l1_in_0_.out ),
    .TE_B(_0159_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.mux_l1_in_1_.out ),
    .TE_B(_0160_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0161_),
    .Z(\cby_0__1_.mux_right_ipin_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_2_.out ),
    .TE_B(_0162_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_3_.out ),
    .TE_B(_0163_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.out ),
    .TE_B(_0164_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_3_.out ),
    .TE_B(_0162_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_4_.out ),
    .TE_B(_0163_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_0164_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_4.mux_l1_in_0_.out ),
    .TE_B(_0165_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_4.mux_l1_in_1_.out ),
    .TE_B(_0166_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0167_),
    .Z(\cby_0__1_.mux_right_ipin_4.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .TE_B(_0168_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0169_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.out ),
    .TE_B(_0170_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_3_.out ),
    .TE_B(_0168_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .TE_B(_0169_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.out ),
    .TE_B(_0170_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_5.mux_l1_in_0_.out ),
    .TE_B(_0171_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_5.mux_l1_in_1_.out ),
    .TE_B(_0172_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0173_),
    .Z(\cby_0__1_.mux_right_ipin_5.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.INVTX1_2_.out ),
    .TE_B(_0174_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.out ),
    .TE_B(_0175_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.INVTX1_4_.out ),
    .TE_B(_0176_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.out ),
    .TE_B(_0174_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_4_.out ),
    .TE_B(_0175_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_5_.out ),
    .TE_B(_0176_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_6.mux_l1_in_0_.out ),
    .TE_B(_0177_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_6.mux_l1_in_1_.out ),
    .TE_B(_0178_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0179_),
    .Z(\cby_0__1_.mux_right_ipin_6.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_2_.out ),
    .TE_B(_0180_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_3_.out ),
    .TE_B(_0181_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_4_.out ),
    .TE_B(_0182_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_0.INVTX1_5_.out ),
    .TE_B(_0180_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0181_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_0__1_.mux_right_ipin_1.INVTX1_5_.out ),
    .TE_B(_0182_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_7.mux_l1_in_0_.out ),
    .TE_B(_0183_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_7.mux_l1_in_1_.out ),
    .TE_B(_0184_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0185_),
    .Z(\cby_0__1_.mux_right_ipin_7.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .TE_B(_0186_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0187_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_2_.out ),
    .TE_B(_0188_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.out ),
    .TE_B(_0186_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_4_.out ),
    .TE_B(_0187_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_0188_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0189_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0190_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0191_),
    .Z(\cby_1__1_.mux_left_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .TE_B(_0192_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0193_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.out ),
    .TE_B(_0194_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0192_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.out ),
    .TE_B(_0193_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_1.INVTX1_5_.out ),
    .TE_B(_0194_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0195_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0196_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0197_),
    .Z(\cby_1__1_.mux_left_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.out ),
    .TE_B(_0198_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0199_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_2_.out ),
    .TE_B(_0200_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0198_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_4_.out ),
    .TE_B(_0199_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_5_.out ),
    .TE_B(_0200_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.mux_l1_in_0_.out ),
    .TE_B(_0201_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.mux_l1_in_1_.out ),
    .TE_B(_0202_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0203_),
    .Z(\cby_1__1_.mux_left_ipin_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_2_.out ),
    .TE_B(_0204_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0205_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_2_.out ),
    .TE_B(_0206_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0204_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_4_.out ),
    .TE_B(_0205_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_5_.out ),
    .TE_B(_0206_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.mux_l1_in_0_.out ),
    .TE_B(_0207_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.mux_l1_in_1_.out ),
    .TE_B(_0208_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0209_),
    .Z(\cby_1__1_.mux_left_ipin_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_2_.out ),
    .TE_B(_0210_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0211_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_2_.out ),
    .TE_B(_0212_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_3_.out ),
    .TE_B(_0210_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_4_.out ),
    .TE_B(_0211_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_5_.out ),
    .TE_B(_0212_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.mux_l1_in_0_.out ),
    .TE_B(_0213_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.mux_l1_in_1_.out ),
    .TE_B(_0214_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0215_),
    .Z(\cby_1__1_.mux_left_ipin_4.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_2_.out ),
    .TE_B(_0216_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_3_.out ),
    .TE_B(_0217_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_2_.out ),
    .TE_B(_0218_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_3_.out ),
    .TE_B(_0216_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_4_.out ),
    .TE_B(_0217_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_5_.out ),
    .TE_B(_0218_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.mux_l1_in_0_.out ),
    .TE_B(_0219_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.mux_l1_in_1_.out ),
    .TE_B(_0220_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0221_),
    .Z(\cby_1__1_.mux_left_ipin_5.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_2_.out ),
    .TE_B(_0222_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_3_.out ),
    .TE_B(_0223_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_2_.out ),
    .TE_B(_0224_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.out ),
    .TE_B(_0222_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_4_.out ),
    .TE_B(_0223_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_0224_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_6.mux_l1_in_0_.out ),
    .TE_B(_0225_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_6.mux_l1_in_1_.out ),
    .TE_B(_0226_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0227_),
    .Z(\cby_1__1_.mux_left_ipin_6.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.out ),
    .TE_B(_0228_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0229_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_2_.out ),
    .TE_B(_0230_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.out ),
    .TE_B(_0228_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.out ),
    .TE_B(_0229_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_1.INVTX1_5_.out ),
    .TE_B(_0230_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_7.mux_l1_in_0_.out ),
    .TE_B(_0231_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_7.mux_l1_in_1_.out ),
    .TE_B(_0232_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0233_),
    .Z(\cby_1__1_.mux_left_ipin_7.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.out ),
    .TE_B(_0234_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0235_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.out ),
    .TE_B(_0236_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_1.INVTX1_5_.out ),
    .TE_B(_0234_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_4_.out ),
    .TE_B(_0235_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_5_.out ),
    .TE_B(_0236_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l1_in_0_.out ),
    .TE_B(_0237_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l1_in_1_.out ),
    .TE_B(_0238_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0239_),
    .Z(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_2_.out ),
    .TE_B(_0240_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0241_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_4_.out ),
    .TE_B(_0242_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_2.INVTX1_5_.out ),
    .TE_B(_0240_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_4_.out ),
    .TE_B(_0241_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_5_.out ),
    .TE_B(_0242_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l1_in_0_.out ),
    .TE_B(_0243_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l1_in_1_.out ),
    .TE_B(_0244_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0245_),
    .Z(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_2_.out ),
    .TE_B(_0246_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0247_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_4_.out ),
    .TE_B(_0248_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_3.INVTX1_5_.out ),
    .TE_B(_0246_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_4_.out ),
    .TE_B(_0247_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cby_1__1_.mux_left_ipin_4.INVTX1_5_.out ),
    .TE_B(_0248_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l1_in_0_.out ),
    .TE_B(_0249_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l1_in_1_.out ),
    .TE_B(_0250_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0251_),
    .Z(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0252_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0253_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0254_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0255_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0256_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0257_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0258_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0259_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0260_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.INVTX1_0_.out ),
    .TE_B(_0261_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.ble4_lut4_0.lut4_0_.lut4_mux_0_.INVTX1_16_.in ),
    .TE_B(_0262_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0263_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0264_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0265_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0266_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0267_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0264_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0265_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0266_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0267_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0264_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0265_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0266_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0267_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0264_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0265_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0266_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_0_.out ),
    .TE_B(_0268_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_1_.out ),
    .TE_B(_0269_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_2_.out ),
    .TE_B(_0270_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l1_in_3_.out ),
    .TE_B(_0271_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_0.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0272_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0273_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0274_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0275_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0272_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0273_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0274_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0275_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0272_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0273_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0274_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0275_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0272_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0273_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0274_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_0_.out ),
    .TE_B(_0276_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_1_.out ),
    .TE_B(_0277_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_2_.out ),
    .TE_B(_0278_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l1_in_3_.out ),
    .TE_B(_0279_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_1.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0280_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0281_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0282_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0283_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0280_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0281_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0282_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0283_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0280_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0281_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0282_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0283_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0280_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0281_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0282_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_0_.out ),
    .TE_B(_0284_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_1_.out ),
    .TE_B(_0285_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_2_.out ),
    .TE_B(_0286_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l1_in_3_.out ),
    .TE_B(_0287_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_2.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0288_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0289_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0290_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0291_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0288_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0289_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0290_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0291_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0288_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0289_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0290_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0291_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0288_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0289_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0290_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_0_.out ),
    .TE_B(_0292_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_1_.out ),
    .TE_B(_0293_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_2_.out ),
    .TE_B(_0294_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l1_in_3_.out ),
    .TE_B(_0295_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_0_in_3.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0296_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0297_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0298_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0299_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0296_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0297_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0298_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0299_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0296_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0297_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0298_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0299_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0296_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0297_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0298_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_0_.out ),
    .TE_B(_0300_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_1_.out ),
    .TE_B(_0301_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_2_.out ),
    .TE_B(_0302_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l1_in_3_.out ),
    .TE_B(_0303_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_0.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0304_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0305_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0306_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0307_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0304_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0305_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0306_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0307_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0304_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0305_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0306_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0307_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0304_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0305_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0306_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_0_.out ),
    .TE_B(_0308_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_1_.out ),
    .TE_B(_0309_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_2_.out ),
    .TE_B(_0310_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l1_in_3_.out ),
    .TE_B(_0311_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_1.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0312_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0313_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0314_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0315_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0312_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0313_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0314_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0315_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0312_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0313_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0314_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0315_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0312_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0313_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0314_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_0_.out ),
    .TE_B(_0316_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_1_.out ),
    .TE_B(_0317_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_2_.out ),
    .TE_B(_0318_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l1_in_3_.out ),
    .TE_B(_0319_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_2.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0320_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0321_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0322_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0323_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0320_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0321_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0322_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0323_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0320_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0321_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0322_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0323_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0320_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0321_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0322_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_0_.out ),
    .TE_B(_0324_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_1_.out ),
    .TE_B(_0325_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_2_.out ),
    .TE_B(_0326_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l1_in_3_.out ),
    .TE_B(_0327_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_1_in_3.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0328_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0329_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0330_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0331_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0328_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0329_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0330_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0331_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0328_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0329_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0330_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0331_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0328_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0329_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0330_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_0_.out ),
    .TE_B(_0332_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_1_.out ),
    .TE_B(_0333_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_2_.out ),
    .TE_B(_0334_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l1_in_3_.out ),
    .TE_B(_0335_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_0.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0336_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0337_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0338_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0339_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0336_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0337_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0338_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0339_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0336_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0337_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0338_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0339_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0336_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0337_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0338_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_0_.out ),
    .TE_B(_0340_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_1_.out ),
    .TE_B(_0341_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_2_.out ),
    .TE_B(_0342_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l1_in_3_.out ),
    .TE_B(_0343_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_1.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0344_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0345_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0346_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0347_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0344_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0345_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0346_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0347_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0344_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0345_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0346_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0347_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0344_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0345_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0346_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_0_.out ),
    .TE_B(_0348_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_1_.out ),
    .TE_B(_0349_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_2_.out ),
    .TE_B(_0350_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l1_in_3_.out ),
    .TE_B(_0351_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_2.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0352_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0353_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0354_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0355_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0352_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0353_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0354_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0355_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0352_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0353_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0354_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0355_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0352_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0353_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0354_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_0_.out ),
    .TE_B(_0356_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_1_.out ),
    .TE_B(_0357_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_2_.out ),
    .TE_B(_0358_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l1_in_3_.out ),
    .TE_B(_0359_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_2_in_3.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0360_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0361_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0362_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0363_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0360_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0361_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0362_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0363_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0360_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0361_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0362_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0363_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0360_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0361_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0362_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_0_.out ),
    .TE_B(_0364_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_1_.out ),
    .TE_B(_0365_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_2_.out ),
    .TE_B(_0366_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l1_in_3_.out ),
    .TE_B(_0367_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_0.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0368_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0369_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0370_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0371_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0368_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0369_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0370_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0371_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0368_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0369_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0370_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0371_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0368_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0369_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0370_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_0_.out ),
    .TE_B(_0372_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_1_.out ),
    .TE_B(_0373_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_2_.out ),
    .TE_B(_0374_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l1_in_3_.out ),
    .TE_B(_0375_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_1.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0376_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0377_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0378_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0379_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0376_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0377_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0378_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0379_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0376_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0377_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0378_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0379_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0376_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0377_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0378_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_0_.out ),
    .TE_B(_0380_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_1_.out ),
    .TE_B(_0381_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_2_.out ),
    .TE_B(_0382_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l1_in_3_.out ),
    .TE_B(_0383_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_2.mux_l2_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0384_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0385_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0386_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.mux_l2_in_0_.out ),
    .TE_B(_0387_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0384_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0385_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0386_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.ebufn  (.A(\cby_0__1_.mux_left_ipin_1.mux_l2_in_0_.out ),
    .TE_B(_0387_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_top_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0384_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.ebufn  (.A(\cby_1__1_.mux_right_ipin_2.mux_l2_in_0_.out ),
    .TE_B(_0385_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0386_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0387_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.TGATE_3_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0384_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0385_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0386_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_0_.out ),
    .TE_B(_0388_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_1_.out ),
    .TE_B(_0389_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_2_.out ),
    .TE_B(_0390_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l1_in_3_.out ),
    .TE_B(_0391_),
    .Z(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.mux_fle_3_in_3.mux_l2_in_0_.TGATE_3_.out ));
 rram_28 rram_wl_0 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[0] ,
    \sb_1__1_.Q_in[13] ,
    \sb_1__1_.Q_in[42] ,
    \cbx_1__1_.Q_in[3] ,
    \cbx_1__1_.Q_in[32] ,
    \cbx_1__1_.Q_in[61] ,
    \sb_0__1_.Q_in[16] ,
    \sb_0__1_.Q_in[45] ,
    \sb_0__0_.Q_in[2] ,
    \sb_0__0_.Q_in[31] ,
    \sb_0__0_.Q_in[60] ,
    \cby_0__1_.Q_in[13] ,
    \cby_0__1_.Q_in[42] ,
    \sb_1__0_.Q_in[3] ,
    \sb_1__0_.Q_in[32] ,
    \sb_1__0_.Q_in[61] ,
    \cbx_1__0_.Q_in[10] ,
    \cbx_1__0_.Q_in[39] ,
    \cby_1__1_.Q_in[2] ,
    \cby_1__1_.Q_in[31] ,
    \cby_1__1_.Q_in[60] ,
    \grid_clb_1__1_.Q_in[23] ,
    \grid_clb_1__1_.Q_in[52] ,
    \grid_clb_1__1_.Q_in[81] ,
    \grid_clb_1__1_.Q_in[110] ,
    \grid_clb_1__1_.Q_in[139] ,
    \grid_clb_1__1_.Q_in[168] ,
    \grid_clb_1__1_.Q_in[197] }));
 rram_28 rram_wl_1 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[1] ,
    \sb_1__1_.Q_in[14] ,
    \sb_1__1_.Q_in[43] ,
    \cbx_1__1_.Q_in[4] ,
    \cbx_1__1_.Q_in[33] ,
    \cbx_1__1_.Q_in[62] ,
    \sb_0__1_.Q_in[17] ,
    \sb_0__1_.Q_in[46] ,
    \sb_0__0_.Q_in[3] ,
    \sb_0__0_.Q_in[32] ,
    \sb_0__0_.Q_in[61] ,
    \cby_0__1_.Q_in[14] ,
    \cby_0__1_.Q_in[43] ,
    \sb_1__0_.Q_in[4] ,
    \sb_1__0_.Q_in[33] ,
    \sb_1__0_.Q_in[62] ,
    \cbx_1__0_.Q_in[11] ,
    \cbx_1__0_.Q_in[40] ,
    \cby_1__1_.Q_in[3] ,
    \cby_1__1_.Q_in[32] ,
    \cby_1__1_.Q_in[61] ,
    \grid_clb_1__1_.Q_in[24] ,
    \grid_clb_1__1_.Q_in[53] ,
    \grid_clb_1__1_.Q_in[82] ,
    \grid_clb_1__1_.Q_in[111] ,
    \grid_clb_1__1_.Q_in[140] ,
    \grid_clb_1__1_.Q_in[169] ,
    \grid_clb_1__1_.Q_in[198] }));
 rram_28 rram_wl_10 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[2] ,
    \sb_1__1_.Q_in[23] ,
    \sb_1__1_.Q_in[52] ,
    \cbx_1__1_.Q_in[13] ,
    \cbx_1__1_.Q_in[42] ,
    \grid_io_top_1__2_.GPIO_DIR[5] ,
    \sb_0__1_.Q_in[26] ,
    \sb_0__1_.Q_in[55] ,
    \sb_0__0_.Q_in[12] ,
    \sb_0__0_.Q_in[41] ,
    \sb_0__0_.Q_in[70] ,
    \cby_0__1_.Q_in[23] ,
    \cby_0__1_.Q_in[52] ,
    \sb_1__0_.Q_in[13] ,
    \sb_1__0_.Q_in[42] ,
    \sb_1__0_.Q_in[71] ,
    \cbx_1__0_.Q_in[20] ,
    \cbx_1__0_.Q_in[49] ,
    \cby_1__1_.Q_in[12] ,
    \cby_1__1_.Q_in[41] ,
    \grid_clb_1__1_.Q_in[4] ,
    \grid_clb_1__1_.Q_in[33] ,
    \grid_clb_1__1_.Q_in[62] ,
    \grid_clb_1__1_.Q_in[91] ,
    \grid_clb_1__1_.Q_in[120] ,
    \grid_clb_1__1_.Q_in[149] ,
    \grid_clb_1__1_.Q_in[178] ,
    \Q27[10] }));
 rram_28 rram_wl_11 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[3] ,
    \sb_1__1_.Q_in[24] ,
    \sb_1__1_.Q_in[53] ,
    \cbx_1__1_.Q_in[14] ,
    \cbx_1__1_.Q_in[43] ,
    \grid_io_top_1__2_.GPIO_DIR[6] ,
    \sb_0__1_.Q_in[27] ,
    \sb_0__1_.Q_in[56] ,
    \sb_0__0_.Q_in[13] ,
    \sb_0__0_.Q_in[42] ,
    \sb_0__0_.Q_in[71] ,
    \cby_0__1_.Q_in[24] ,
    \cby_0__1_.Q_in[53] ,
    \sb_1__0_.Q_in[14] ,
    \sb_1__0_.Q_in[43] ,
    \sb_1__0_.Q_in[72] ,
    \cbx_1__0_.Q_in[21] ,
    \cbx_1__0_.Q_in[50] ,
    \cby_1__1_.Q_in[13] ,
    \cby_1__1_.Q_in[42] ,
    \grid_clb_1__1_.Q_in[5] ,
    \grid_clb_1__1_.Q_in[34] ,
    \grid_clb_1__1_.Q_in[63] ,
    \grid_clb_1__1_.Q_in[92] ,
    \grid_clb_1__1_.Q_in[121] ,
    \grid_clb_1__1_.Q_in[150] ,
    \grid_clb_1__1_.Q_in[179] ,
    \Q27[11] }));
 rram_28 rram_wl_12 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[4] ,
    \sb_1__1_.Q_in[25] ,
    \sb_1__1_.Q_in[54] ,
    \cbx_1__1_.Q_in[15] ,
    \cbx_1__1_.Q_in[44] ,
    \grid_io_top_1__2_.GPIO_DIR[7] ,
    \sb_0__1_.Q_in[28] ,
    \sb_0__1_.Q_in[57] ,
    \sb_0__0_.Q_in[14] ,
    \sb_0__0_.Q_in[43] ,
    \sb_0__0_.Q_in[72] ,
    \cby_0__1_.Q_in[25] ,
    \cby_0__1_.Q_in[54] ,
    \sb_1__0_.Q_in[15] ,
    \sb_1__0_.Q_in[44] ,
    \sb_1__0_.Q_in[73] ,
    \cbx_1__0_.Q_in[22] ,
    \cbx_1__0_.Q_in[51] ,
    \cby_1__1_.Q_in[14] ,
    \cby_1__1_.Q_in[43] ,
    \grid_clb_1__1_.Q_in[6] ,
    \grid_clb_1__1_.Q_in[35] ,
    \grid_clb_1__1_.Q_in[64] ,
    \grid_clb_1__1_.Q_in[93] ,
    \grid_clb_1__1_.Q_in[122] ,
    \grid_clb_1__1_.Q_in[151] ,
    \grid_clb_1__1_.Q_in[180] ,
    \Q27[12] }));
 rram_28 rram_wl_13 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[5] ,
    \sb_1__1_.Q_in[26] ,
    \sb_1__1_.Q_in[55] ,
    \cbx_1__1_.Q_in[16] ,
    \cbx_1__1_.Q_in[45] ,
    \Q5[13] ,
    \sb_0__1_.Q_in[29] ,
    \sb_0__1_.Q_in[58] ,
    \sb_0__0_.Q_in[15] ,
    \sb_0__0_.Q_in[44] ,
    \sb_0__0_.Q_in[73] ,
    \cby_0__1_.Q_in[26] ,
    \cby_0__1_.Q_in[55] ,
    \sb_1__0_.Q_in[16] ,
    \sb_1__0_.Q_in[45] ,
    \sb_1__0_.Q_in[74] ,
    \cbx_1__0_.Q_in[23] ,
    \cbx_1__0_.Q_in[52] ,
    \cby_1__1_.Q_in[15] ,
    \cby_1__1_.Q_in[44] ,
    \grid_clb_1__1_.Q_in[7] ,
    \grid_clb_1__1_.Q_in[36] ,
    \grid_clb_1__1_.Q_in[65] ,
    \grid_clb_1__1_.Q_in[94] ,
    \grid_clb_1__1_.Q_in[123] ,
    \grid_clb_1__1_.Q_in[152] ,
    \grid_clb_1__1_.Q_in[181] ,
    \Q27[13] }));
 rram_28 rram_wl_14 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[6] ,
    \sb_1__1_.Q_in[27] ,
    \sb_1__1_.Q_in[56] ,
    \cbx_1__1_.Q_in[17] ,
    \cbx_1__1_.Q_in[46] ,
    \Q5[14] ,
    \sb_0__1_.Q_in[30] ,
    \sb_0__1_.Q_in[59] ,
    \sb_0__0_.Q_in[16] ,
    \sb_0__0_.Q_in[45] ,
    \sb_0__0_.Q_in[74] ,
    \cby_0__1_.Q_in[27] ,
    \cby_0__1_.Q_in[56] ,
    \sb_1__0_.Q_in[17] ,
    \sb_1__0_.Q_in[46] ,
    \sb_1__0_.Q_in[75] ,
    \cbx_1__0_.Q_in[24] ,
    \cbx_1__0_.Q_in[53] ,
    \cby_1__1_.Q_in[16] ,
    \cby_1__1_.Q_in[45] ,
    \grid_clb_1__1_.Q_in[8] ,
    \grid_clb_1__1_.Q_in[37] ,
    \grid_clb_1__1_.Q_in[66] ,
    \grid_clb_1__1_.Q_in[95] ,
    \grid_clb_1__1_.Q_in[124] ,
    \grid_clb_1__1_.Q_in[153] ,
    \grid_clb_1__1_.Q_in[182] ,
    \Q27[14] }));
 rram_28 rram_wl_15 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[7] ,
    \sb_1__1_.Q_in[28] ,
    \sb_1__1_.Q_in[57] ,
    \cbx_1__1_.Q_in[18] ,
    \cbx_1__1_.Q_in[47] ,
    \Q5[15] ,
    \sb_0__1_.Q_in[31] ,
    \sb_0__1_.Q_in[60] ,
    \sb_0__0_.Q_in[17] ,
    \sb_0__0_.Q_in[46] ,
    \sb_0__0_.Q_in[75] ,
    \cby_0__1_.Q_in[28] ,
    \cby_0__1_.Q_in[57] ,
    \sb_1__0_.Q_in[18] ,
    \sb_1__0_.Q_in[47] ,
    \sb_1__0_.Q_in[76] ,
    \cbx_1__0_.Q_in[25] ,
    \cbx_1__0_.Q_in[54] ,
    \cby_1__1_.Q_in[17] ,
    \cby_1__1_.Q_in[46] ,
    \grid_clb_1__1_.Q_in[9] ,
    \grid_clb_1__1_.Q_in[38] ,
    \grid_clb_1__1_.Q_in[67] ,
    \grid_clb_1__1_.Q_in[96] ,
    \grid_clb_1__1_.Q_in[125] ,
    \grid_clb_1__1_.Q_in[154] ,
    \grid_clb_1__1_.Q_in[183] ,
    \Q27[15] }));
 rram_28 rram_wl_16 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[0] ,
    \sb_1__1_.Q_in[29] ,
    \sb_1__1_.Q_in[58] ,
    \cbx_1__1_.Q_in[19] ,
    \cbx_1__1_.Q_in[48] ,
    \Q5[16] ,
    \sb_0__1_.Q_in[32] ,
    \sb_0__1_.Q_in[61] ,
    \sb_0__0_.Q_in[18] ,
    \sb_0__0_.Q_in[47] ,
    \cby_0__1_.Q_in[0] ,
    \cby_0__1_.Q_in[29] ,
    \cby_0__1_.Q_in[58] ,
    \sb_1__0_.Q_in[19] ,
    \sb_1__0_.Q_in[48] ,
    \sb_1__0_.Q_in[77] ,
    \cbx_1__0_.Q_in[26] ,
    \cbx_1__0_.Q_in[55] ,
    \cby_1__1_.Q_in[18] ,
    \cby_1__1_.Q_in[47] ,
    \grid_clb_1__1_.Q_in[10] ,
    \grid_clb_1__1_.Q_in[39] ,
    \grid_clb_1__1_.Q_in[68] ,
    \grid_clb_1__1_.Q_in[97] ,
    \grid_clb_1__1_.Q_in[126] ,
    \grid_clb_1__1_.Q_in[155] ,
    \grid_clb_1__1_.Q_in[184] ,
    \Q27[16] }));
 rram_28 rram_wl_17 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[1] ,
    \sb_1__1_.Q_in[30] ,
    \sb_1__1_.Q_in[59] ,
    \cbx_1__1_.Q_in[20] ,
    \cbx_1__1_.Q_in[49] ,
    \Q5[17] ,
    \sb_0__1_.Q_in[33] ,
    \sb_0__1_.Q_in[62] ,
    \sb_0__0_.Q_in[19] ,
    \sb_0__0_.Q_in[48] ,
    \cby_0__1_.Q_in[1] ,
    \cby_0__1_.Q_in[30] ,
    \cby_0__1_.Q_in[59] ,
    \sb_1__0_.Q_in[20] ,
    \sb_1__0_.Q_in[49] ,
    \sb_1__0_.Q_in[78] ,
    \cbx_1__0_.Q_in[27] ,
    \cbx_1__0_.Q_in[56] ,
    \cby_1__1_.Q_in[19] ,
    \cby_1__1_.Q_in[48] ,
    \grid_clb_1__1_.Q_in[11] ,
    \grid_clb_1__1_.Q_in[40] ,
    \grid_clb_1__1_.Q_in[69] ,
    \grid_clb_1__1_.Q_in[98] ,
    \grid_clb_1__1_.Q_in[127] ,
    \grid_clb_1__1_.Q_in[156] ,
    \grid_clb_1__1_.Q_in[185] ,
    \Q27[17] }));
 rram_28 rram_wl_18 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[2] ,
    \sb_1__1_.Q_in[31] ,
    \sb_1__1_.Q_in[60] ,
    \cbx_1__1_.Q_in[21] ,
    \cbx_1__1_.Q_in[50] ,
    \Q5[18] ,
    \sb_0__1_.Q_in[34] ,
    \sb_0__1_.Q_in[63] ,
    \sb_0__0_.Q_in[20] ,
    \sb_0__0_.Q_in[49] ,
    \cby_0__1_.Q_in[2] ,
    \cby_0__1_.Q_in[31] ,
    \grid_io_left_0__1_.GPIO_DIR[0] ,
    \sb_1__0_.Q_in[21] ,
    \sb_1__0_.Q_in[50] ,
    \sb_1__0_.Q_in[79] ,
    \cbx_1__0_.Q_in[28] ,
    \cbx_1__0_.Q_in[57] ,
    \cby_1__1_.Q_in[20] ,
    \cby_1__1_.Q_in[49] ,
    \grid_clb_1__1_.Q_in[12] ,
    \grid_clb_1__1_.Q_in[41] ,
    \grid_clb_1__1_.Q_in[70] ,
    \grid_clb_1__1_.Q_in[99] ,
    \grid_clb_1__1_.Q_in[128] ,
    \grid_clb_1__1_.Q_in[157] ,
    \grid_clb_1__1_.Q_in[186] ,
    \Q27[18] }));
 rram_28 rram_wl_19 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[3] ,
    \sb_1__1_.Q_in[32] ,
    \sb_1__1_.Q_in[61] ,
    \cbx_1__1_.Q_in[22] ,
    \cbx_1__1_.Q_in[51] ,
    \Q5[19] ,
    \sb_0__1_.Q_in[35] ,
    \sb_0__1_.Q_in[64] ,
    \sb_0__0_.Q_in[21] ,
    \sb_0__0_.Q_in[50] ,
    \cby_0__1_.Q_in[3] ,
    \cby_0__1_.Q_in[32] ,
    \grid_io_left_0__1_.GPIO_DIR[1] ,
    \sb_1__0_.Q_in[22] ,
    \sb_1__0_.Q_in[51] ,
    \cbx_1__0_.Q_in[0] ,
    \cbx_1__0_.Q_in[29] ,
    \cbx_1__0_.Q_in[58] ,
    \cby_1__1_.Q_in[21] ,
    \cby_1__1_.Q_in[50] ,
    \grid_clb_1__1_.Q_in[13] ,
    \grid_clb_1__1_.Q_in[42] ,
    \grid_clb_1__1_.Q_in[71] ,
    \grid_clb_1__1_.Q_in[100] ,
    \grid_clb_1__1_.Q_in[129] ,
    \grid_clb_1__1_.Q_in[158] ,
    \grid_clb_1__1_.Q_in[187] ,
    \Q27[19] }));
 rram_28 rram_wl_2 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[2] ,
    \sb_1__1_.Q_in[15] ,
    \sb_1__1_.Q_in[44] ,
    \cbx_1__1_.Q_in[5] ,
    \cbx_1__1_.Q_in[34] ,
    \cbx_1__1_.Q_in[63] ,
    \sb_0__1_.Q_in[18] ,
    \sb_0__1_.Q_in[47] ,
    \sb_0__0_.Q_in[4] ,
    \sb_0__0_.Q_in[33] ,
    \sb_0__0_.Q_in[62] ,
    \cby_0__1_.Q_in[15] ,
    \cby_0__1_.Q_in[44] ,
    \sb_1__0_.Q_in[5] ,
    \sb_1__0_.Q_in[34] ,
    \sb_1__0_.Q_in[63] ,
    \cbx_1__0_.Q_in[12] ,
    \cbx_1__0_.Q_in[41] ,
    \cby_1__1_.Q_in[4] ,
    \cby_1__1_.Q_in[33] ,
    \cby_1__1_.Q_in[62] ,
    \grid_clb_1__1_.Q_in[25] ,
    \grid_clb_1__1_.Q_in[54] ,
    \grid_clb_1__1_.Q_in[83] ,
    \grid_clb_1__1_.Q_in[112] ,
    \grid_clb_1__1_.Q_in[141] ,
    \grid_clb_1__1_.Q_in[170] ,
    \grid_clb_1__1_.Q_in[199] }));
 rram_28 rram_wl_20 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[4] ,
    \sb_1__1_.Q_in[33] ,
    \sb_1__1_.Q_in[62] ,
    \cbx_1__1_.Q_in[23] ,
    \cbx_1__1_.Q_in[52] ,
    \Q5[20] ,
    \sb_0__1_.Q_in[36] ,
    \sb_0__1_.Q_in[65] ,
    \sb_0__0_.Q_in[22] ,
    \sb_0__0_.Q_in[51] ,
    \cby_0__1_.Q_in[4] ,
    \cby_0__1_.Q_in[33] ,
    \grid_io_left_0__1_.GPIO_DIR[2] ,
    \sb_1__0_.Q_in[23] ,
    \sb_1__0_.Q_in[52] ,
    \cbx_1__0_.Q_in[1] ,
    \cbx_1__0_.Q_in[30] ,
    \cbx_1__0_.Q_in[59] ,
    \cby_1__1_.Q_in[22] ,
    \cby_1__1_.Q_in[51] ,
    \grid_clb_1__1_.Q_in[14] ,
    \grid_clb_1__1_.Q_in[43] ,
    \grid_clb_1__1_.Q_in[72] ,
    \grid_clb_1__1_.Q_in[101] ,
    \grid_clb_1__1_.Q_in[130] ,
    \grid_clb_1__1_.Q_in[159] ,
    \grid_clb_1__1_.Q_in[188] ,
    \Q27[20] }));
 rram_28 rram_wl_21 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[5] ,
    \sb_1__1_.Q_in[34] ,
    \sb_1__1_.Q_in[63] ,
    \cbx_1__1_.Q_in[24] ,
    \cbx_1__1_.Q_in[53] ,
    \Q5[21] ,
    \sb_0__1_.Q_in[37] ,
    \sb_0__1_.Q_in[66] ,
    \sb_0__0_.Q_in[23] ,
    \sb_0__0_.Q_in[52] ,
    \cby_0__1_.Q_in[5] ,
    \cby_0__1_.Q_in[34] ,
    \grid_io_left_0__1_.GPIO_DIR[3] ,
    \sb_1__0_.Q_in[24] ,
    \sb_1__0_.Q_in[53] ,
    \cbx_1__0_.Q_in[2] ,
    \cbx_1__0_.Q_in[31] ,
    \cbx_1__0_.Q_in[60] ,
    \cby_1__1_.Q_in[23] ,
    \cby_1__1_.Q_in[52] ,
    \grid_clb_1__1_.Q_in[15] ,
    \grid_clb_1__1_.Q_in[44] ,
    \grid_clb_1__1_.Q_in[73] ,
    \grid_clb_1__1_.Q_in[102] ,
    \grid_clb_1__1_.Q_in[131] ,
    \grid_clb_1__1_.Q_in[160] ,
    \grid_clb_1__1_.Q_in[189] ,
    \Q27[21] }));
 rram_28 rram_wl_22 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[6] ,
    \sb_1__1_.Q_in[35] ,
    \sb_1__1_.Q_in[64] ,
    \cbx_1__1_.Q_in[25] ,
    \cbx_1__1_.Q_in[54] ,
    \Q5[22] ,
    \sb_0__1_.Q_in[38] ,
    \sb_0__1_.Q_in[67] ,
    \sb_0__0_.Q_in[24] ,
    \sb_0__0_.Q_in[53] ,
    \cby_0__1_.Q_in[6] ,
    \cby_0__1_.Q_in[35] ,
    \grid_io_left_0__1_.GPIO_DIR[4] ,
    \sb_1__0_.Q_in[25] ,
    \sb_1__0_.Q_in[54] ,
    \cbx_1__0_.Q_in[3] ,
    \cbx_1__0_.Q_in[32] ,
    \cbx_1__0_.Q_in[61] ,
    \cby_1__1_.Q_in[24] ,
    \cby_1__1_.Q_in[53] ,
    \grid_clb_1__1_.Q_in[16] ,
    \grid_clb_1__1_.Q_in[45] ,
    \grid_clb_1__1_.Q_in[74] ,
    \grid_clb_1__1_.Q_in[103] ,
    \grid_clb_1__1_.Q_in[132] ,
    \grid_clb_1__1_.Q_in[161] ,
    \grid_clb_1__1_.Q_in[190] ,
    \Q27[22] }));
 rram_28 rram_wl_23 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[7] ,
    \sb_1__1_.Q_in[36] ,
    \sb_1__1_.Q_in[65] ,
    \cbx_1__1_.Q_in[26] ,
    \cbx_1__1_.Q_in[55] ,
    \Q5[23] ,
    \sb_0__1_.Q_in[39] ,
    \sb_0__1_.Q_in[68] ,
    \sb_0__0_.Q_in[25] ,
    \sb_0__0_.Q_in[54] ,
    \cby_0__1_.Q_in[7] ,
    \cby_0__1_.Q_in[36] ,
    \grid_io_left_0__1_.GPIO_DIR[5] ,
    \sb_1__0_.Q_in[26] ,
    \sb_1__0_.Q_in[55] ,
    \cbx_1__0_.Q_in[4] ,
    \cbx_1__0_.Q_in[33] ,
    \cbx_1__0_.Q_in[62] ,
    \cby_1__1_.Q_in[25] ,
    \cby_1__1_.Q_in[54] ,
    \grid_clb_1__1_.Q_in[17] ,
    \grid_clb_1__1_.Q_in[46] ,
    \grid_clb_1__1_.Q_in[75] ,
    \grid_clb_1__1_.Q_in[104] ,
    \grid_clb_1__1_.Q_in[133] ,
    \grid_clb_1__1_.Q_in[162] ,
    \grid_clb_1__1_.Q_in[191] ,
    \Q27[23] }));
 rram_28 rram_wl_24 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[8] ,
    \sb_1__1_.Q_in[37] ,
    \sb_1__1_.Q_in[66] ,
    \cbx_1__1_.Q_in[27] ,
    \cbx_1__1_.Q_in[56] ,
    \Q5[24] ,
    \sb_0__1_.Q_in[40] ,
    \sb_0__1_.Q_in[69] ,
    \sb_0__0_.Q_in[26] ,
    \sb_0__0_.Q_in[55] ,
    \cby_0__1_.Q_in[8] ,
    \cby_0__1_.Q_in[37] ,
    \grid_io_left_0__1_.GPIO_DIR[6] ,
    \sb_1__0_.Q_in[27] ,
    \sb_1__0_.Q_in[56] ,
    \cbx_1__0_.Q_in[5] ,
    \cbx_1__0_.Q_in[34] ,
    \cbx_1__0_.Q_in[63] ,
    \cby_1__1_.Q_in[26] ,
    \cby_1__1_.Q_in[55] ,
    \grid_clb_1__1_.Q_in[18] ,
    \grid_clb_1__1_.Q_in[47] ,
    \grid_clb_1__1_.Q_in[76] ,
    \grid_clb_1__1_.Q_in[105] ,
    \grid_clb_1__1_.Q_in[134] ,
    \grid_clb_1__1_.Q_in[163] ,
    \grid_clb_1__1_.Q_in[192] ,
    \Q27[24] }));
 rram_28 rram_wl_25 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[9] ,
    \sb_1__1_.Q_in[38] ,
    \sb_1__1_.Q_in[67] ,
    \cbx_1__1_.Q_in[28] ,
    \cbx_1__1_.Q_in[57] ,
    \Q5[25] ,
    \sb_0__1_.Q_in[41] ,
    \sb_0__1_.Q_in[70] ,
    \sb_0__0_.Q_in[27] ,
    \sb_0__0_.Q_in[56] ,
    \cby_0__1_.Q_in[9] ,
    \cby_0__1_.Q_in[38] ,
    \grid_io_left_0__1_.GPIO_DIR[7] ,
    \sb_1__0_.Q_in[28] ,
    \sb_1__0_.Q_in[57] ,
    \cbx_1__0_.Q_in[6] ,
    \cbx_1__0_.Q_in[35] ,
    \cbx_1__0_.Q_in[64] ,
    \cby_1__1_.Q_in[27] ,
    \cby_1__1_.Q_in[56] ,
    \grid_clb_1__1_.Q_in[19] ,
    \grid_clb_1__1_.Q_in[48] ,
    \grid_clb_1__1_.Q_in[77] ,
    \grid_clb_1__1_.Q_in[106] ,
    \grid_clb_1__1_.Q_in[135] ,
    \grid_clb_1__1_.Q_in[164] ,
    \grid_clb_1__1_.Q_in[193] ,
    \Q27[25] }));
 rram_28 rram_wl_26 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[10] ,
    \sb_1__1_.Q_in[39] ,
    \cbx_1__1_.Q_in[0] ,
    \cbx_1__1_.Q_in[29] ,
    \cbx_1__1_.Q_in[58] ,
    \Q5[26] ,
    \sb_0__1_.Q_in[42] ,
    \sb_0__1_.Q_in[71] ,
    \sb_0__0_.Q_in[28] ,
    \sb_0__0_.Q_in[57] ,
    \cby_0__1_.Q_in[10] ,
    \cby_0__1_.Q_in[39] ,
    \sb_1__0_.Q_in[0] ,
    \sb_1__0_.Q_in[29] ,
    \sb_1__0_.Q_in[58] ,
    \cbx_1__0_.Q_in[7] ,
    \cbx_1__0_.Q_in[36] ,
    \cbx_1__0_.Q_in[65] ,
    \cby_1__1_.Q_in[28] ,
    \cby_1__1_.Q_in[57] ,
    \grid_clb_1__1_.Q_in[20] ,
    \grid_clb_1__1_.Q_in[49] ,
    \grid_clb_1__1_.Q_in[78] ,
    \grid_clb_1__1_.Q_in[107] ,
    \grid_clb_1__1_.Q_in[136] ,
    \grid_clb_1__1_.Q_in[165] ,
    \grid_clb_1__1_.Q_in[194] ,
    \Q27[26] }));
 rram_28 rram_wl_27 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[11] ,
    \sb_1__1_.Q_in[40] ,
    \cbx_1__1_.Q_in[1] ,
    \cbx_1__1_.Q_in[30] ,
    \cbx_1__1_.Q_in[59] ,
    \sb_0__1_.Q_in[14] ,
    \sb_0__1_.Q_in[43] ,
    \sb_0__0_.Q_in[0] ,
    \sb_0__0_.Q_in[29] ,
    \sb_0__0_.Q_in[58] ,
    \cby_0__1_.Q_in[11] ,
    \cby_0__1_.Q_in[40] ,
    \sb_1__0_.Q_in[1] ,
    \sb_1__0_.Q_in[30] ,
    \sb_1__0_.Q_in[59] ,
    \cbx_1__0_.Q_in[8] ,
    \cbx_1__0_.Q_in[37] ,
    \cby_1__1_.Q_in[0] ,
    \cby_1__1_.Q_in[29] ,
    \cby_1__1_.Q_in[58] ,
    \grid_clb_1__1_.Q_in[21] ,
    \grid_clb_1__1_.Q_in[50] ,
    \grid_clb_1__1_.Q_in[79] ,
    \grid_clb_1__1_.Q_in[108] ,
    \grid_clb_1__1_.Q_in[137] ,
    \grid_clb_1__1_.Q_in[166] ,
    \grid_clb_1__1_.Q_in[195] ,
    \Q27[27] }));
 rram_28 rram_wl_28 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\sb_1__1_.Q_in[12] ,
    \sb_1__1_.Q_in[41] ,
    \cbx_1__1_.Q_in[2] ,
    \cbx_1__1_.Q_in[31] ,
    \cbx_1__1_.Q_in[60] ,
    \sb_0__1_.Q_in[15] ,
    \sb_0__1_.Q_in[44] ,
    \sb_0__0_.Q_in[1] ,
    \sb_0__0_.Q_in[30] ,
    \sb_0__0_.Q_in[59] ,
    \cby_0__1_.Q_in[12] ,
    \cby_0__1_.Q_in[41] ,
    \sb_1__0_.Q_in[2] ,
    \sb_1__0_.Q_in[31] ,
    \sb_1__0_.Q_in[60] ,
    \cbx_1__0_.Q_in[9] ,
    \cbx_1__0_.Q_in[38] ,
    \cby_1__1_.Q_in[1] ,
    \cby_1__1_.Q_in[30] ,
    \cby_1__1_.Q_in[59] ,
    \grid_clb_1__1_.Q_in[22] ,
    \grid_clb_1__1_.Q_in[51] ,
    \grid_clb_1__1_.Q_in[80] ,
    \grid_clb_1__1_.Q_in[109] ,
    \grid_clb_1__1_.Q_in[138] ,
    \grid_clb_1__1_.Q_in[167] ,
    \grid_clb_1__1_.Q_in[196] ,
    \Q27[28] }));
 rram_28 rram_wl_3 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[3] ,
    \sb_1__1_.Q_in[16] ,
    \sb_1__1_.Q_in[45] ,
    \cbx_1__1_.Q_in[6] ,
    \cbx_1__1_.Q_in[35] ,
    \cbx_1__1_.Q_in[64] ,
    \sb_0__1_.Q_in[19] ,
    \sb_0__1_.Q_in[48] ,
    \sb_0__0_.Q_in[5] ,
    \sb_0__0_.Q_in[34] ,
    \sb_0__0_.Q_in[63] ,
    \cby_0__1_.Q_in[16] ,
    \cby_0__1_.Q_in[45] ,
    \sb_1__0_.Q_in[6] ,
    \sb_1__0_.Q_in[35] ,
    \sb_1__0_.Q_in[64] ,
    \cbx_1__0_.Q_in[13] ,
    \cbx_1__0_.Q_in[42] ,
    \cby_1__1_.Q_in[5] ,
    \cby_1__1_.Q_in[34] ,
    \cby_1__1_.Q_in[63] ,
    \grid_clb_1__1_.Q_in[26] ,
    \grid_clb_1__1_.Q_in[55] ,
    \grid_clb_1__1_.Q_in[84] ,
    \grid_clb_1__1_.Q_in[113] ,
    \grid_clb_1__1_.Q_in[142] ,
    \grid_clb_1__1_.Q_in[171] ,
    \grid_clb_1__1_.Q_in[200] }));
 rram_28 rram_wl_4 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[4] ,
    \sb_1__1_.Q_in[17] ,
    \sb_1__1_.Q_in[46] ,
    \cbx_1__1_.Q_in[7] ,
    \cbx_1__1_.Q_in[36] ,
    \cbx_1__1_.Q_in[65] ,
    \sb_0__1_.Q_in[20] ,
    \sb_0__1_.Q_in[49] ,
    \sb_0__0_.Q_in[6] ,
    \sb_0__0_.Q_in[35] ,
    \sb_0__0_.Q_in[64] ,
    \cby_0__1_.Q_in[17] ,
    \cby_0__1_.Q_in[46] ,
    \sb_1__0_.Q_in[7] ,
    \sb_1__0_.Q_in[36] ,
    \sb_1__0_.Q_in[65] ,
    \cbx_1__0_.Q_in[14] ,
    \cbx_1__0_.Q_in[43] ,
    \cby_1__1_.Q_in[6] ,
    \cby_1__1_.Q_in[35] ,
    \cby_1__1_.Q_in[64] ,
    \grid_clb_1__1_.Q_in[27] ,
    \grid_clb_1__1_.Q_in[56] ,
    \grid_clb_1__1_.Q_in[85] ,
    \grid_clb_1__1_.Q_in[114] ,
    \grid_clb_1__1_.Q_in[143] ,
    \grid_clb_1__1_.Q_in[172] ,
    \grid_clb_1__1_.Q_in[201] }));
 rram_28 rram_wl_5 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[5] ,
    \sb_1__1_.Q_in[18] ,
    \sb_1__1_.Q_in[47] ,
    \cbx_1__1_.Q_in[8] ,
    \cbx_1__1_.Q_in[37] ,
    \grid_io_top_1__2_.GPIO_DIR[0] ,
    \sb_0__1_.Q_in[21] ,
    \sb_0__1_.Q_in[50] ,
    \sb_0__0_.Q_in[7] ,
    \sb_0__0_.Q_in[36] ,
    \sb_0__0_.Q_in[65] ,
    \cby_0__1_.Q_in[18] ,
    \cby_0__1_.Q_in[47] ,
    \sb_1__0_.Q_in[8] ,
    \sb_1__0_.Q_in[37] ,
    \sb_1__0_.Q_in[66] ,
    \cbx_1__0_.Q_in[15] ,
    \cbx_1__0_.Q_in[44] ,
    \cby_1__1_.Q_in[7] ,
    \cby_1__1_.Q_in[36] ,
    \cby_1__1_.Q_in[65] ,
    \grid_clb_1__1_.Q_in[28] ,
    \grid_clb_1__1_.Q_in[57] ,
    \grid_clb_1__1_.Q_in[86] ,
    \grid_clb_1__1_.Q_in[115] ,
    \grid_clb_1__1_.Q_in[144] ,
    \grid_clb_1__1_.Q_in[173] ,
    \grid_clb_1__1_.Q_in[202] }));
 rram_28 rram_wl_6 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[6] ,
    \sb_1__1_.Q_in[19] ,
    \sb_1__1_.Q_in[48] ,
    \cbx_1__1_.Q_in[9] ,
    \cbx_1__1_.Q_in[38] ,
    \grid_io_top_1__2_.GPIO_DIR[1] ,
    \sb_0__1_.Q_in[22] ,
    \sb_0__1_.Q_in[51] ,
    \sb_0__0_.Q_in[8] ,
    \sb_0__0_.Q_in[37] ,
    \sb_0__0_.Q_in[66] ,
    \cby_0__1_.Q_in[19] ,
    \cby_0__1_.Q_in[48] ,
    \sb_1__0_.Q_in[9] ,
    \sb_1__0_.Q_in[38] ,
    \sb_1__0_.Q_in[67] ,
    \cbx_1__0_.Q_in[16] ,
    \cbx_1__0_.Q_in[45] ,
    \cby_1__1_.Q_in[8] ,
    \cby_1__1_.Q_in[37] ,
    \grid_clb_1__1_.Q_in[0] ,
    \grid_clb_1__1_.Q_in[29] ,
    \grid_clb_1__1_.Q_in[58] ,
    \grid_clb_1__1_.Q_in[87] ,
    \grid_clb_1__1_.Q_in[116] ,
    \grid_clb_1__1_.Q_in[145] ,
    \grid_clb_1__1_.Q_in[174] ,
    \grid_clb_1__1_.Q_in[203] }));
 rram_28 rram_wl_7 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_bottom_1__0_.GPIO_DIR[7] ,
    \sb_1__1_.Q_in[20] ,
    \sb_1__1_.Q_in[49] ,
    \cbx_1__1_.Q_in[10] ,
    \cbx_1__1_.Q_in[39] ,
    \grid_io_top_1__2_.GPIO_DIR[2] ,
    \sb_0__1_.Q_in[23] ,
    \sb_0__1_.Q_in[52] ,
    \sb_0__0_.Q_in[9] ,
    \sb_0__0_.Q_in[38] ,
    \sb_0__0_.Q_in[67] ,
    \cby_0__1_.Q_in[20] ,
    \cby_0__1_.Q_in[49] ,
    \sb_1__0_.Q_in[10] ,
    \sb_1__0_.Q_in[39] ,
    \sb_1__0_.Q_in[68] ,
    \cbx_1__0_.Q_in[17] ,
    \cbx_1__0_.Q_in[46] ,
    \cby_1__1_.Q_in[9] ,
    \cby_1__1_.Q_in[38] ,
    \grid_clb_1__1_.Q_in[1] ,
    \grid_clb_1__1_.Q_in[30] ,
    \grid_clb_1__1_.Q_in[59] ,
    \grid_clb_1__1_.Q_in[88] ,
    \grid_clb_1__1_.Q_in[117] ,
    \grid_clb_1__1_.Q_in[146] ,
    \grid_clb_1__1_.Q_in[175] ,
    \Q27[7] }));
 rram_28 rram_wl_8 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[0] ,
    \sb_1__1_.Q_in[21] ,
    \sb_1__1_.Q_in[50] ,
    \cbx_1__1_.Q_in[11] ,
    \cbx_1__1_.Q_in[40] ,
    \grid_io_top_1__2_.GPIO_DIR[3] ,
    \sb_0__1_.Q_in[24] ,
    \sb_0__1_.Q_in[53] ,
    \sb_0__0_.Q_in[10] ,
    \sb_0__0_.Q_in[39] ,
    \sb_0__0_.Q_in[68] ,
    \cby_0__1_.Q_in[21] ,
    \cby_0__1_.Q_in[50] ,
    \sb_1__0_.Q_in[11] ,
    \sb_1__0_.Q_in[40] ,
    \sb_1__0_.Q_in[69] ,
    \cbx_1__0_.Q_in[18] ,
    \cbx_1__0_.Q_in[47] ,
    \cby_1__1_.Q_in[10] ,
    \cby_1__1_.Q_in[39] ,
    \grid_clb_1__1_.Q_in[2] ,
    \grid_clb_1__1_.Q_in[31] ,
    \grid_clb_1__1_.Q_in[60] ,
    \grid_clb_1__1_.Q_in[89] ,
    \grid_clb_1__1_.Q_in[118] ,
    \grid_clb_1__1_.Q_in[147] ,
    \grid_clb_1__1_.Q_in[176] ,
    \Q27[8] }));
 rram_28 rram_wl_9 (.BL({data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in,
    data_in}),
    .Q({\grid_io_right_2__1_.GPIO_DIR[1] ,
    \sb_1__1_.Q_in[22] ,
    \sb_1__1_.Q_in[51] ,
    \cbx_1__1_.Q_in[12] ,
    \cbx_1__1_.Q_in[41] ,
    \grid_io_top_1__2_.GPIO_DIR[4] ,
    \sb_0__1_.Q_in[25] ,
    \sb_0__1_.Q_in[54] ,
    \sb_0__0_.Q_in[11] ,
    \sb_0__0_.Q_in[40] ,
    \sb_0__0_.Q_in[69] ,
    \cby_0__1_.Q_in[22] ,
    \cby_0__1_.Q_in[51] ,
    \sb_1__0_.Q_in[12] ,
    \sb_1__0_.Q_in[41] ,
    \sb_1__0_.Q_in[70] ,
    \cbx_1__0_.Q_in[19] ,
    \cbx_1__0_.Q_in[48] ,
    \cby_1__1_.Q_in[11] ,
    \cby_1__1_.Q_in[40] ,
    \grid_clb_1__1_.Q_in[3] ,
    \grid_clb_1__1_.Q_in[32] ,
    \grid_clb_1__1_.Q_in[61] ,
    \grid_clb_1__1_.Q_in[90] ,
    \grid_clb_1__1_.Q_in[119] ,
    \grid_clb_1__1_.Q_in[148] ,
    \grid_clb_1__1_.Q_in[177] ,
    \Q27[9] }));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_0392_),
    .Z(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0393_),
    .Z(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0394_),
    .Z(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_0.mux_l1_in_0_.out ),
    .TE_B(_0395_),
    .Z(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0396_),
    .Z(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0397_),
    .Z(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_3_.out ),
    .TE_B(_0398_),
    .Z(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0399_),
    .Z(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0400_),
    .Z(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_12.mux_l1_in_0_.out ),
    .TE_B(_0401_),
    .Z(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0402_),
    .Z(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0403_),
    .Z(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_0__1_.mux_left_ipin_0.INVTX1_3_.out ),
    .TE_B(_0404_),
    .Z(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0405_),
    .Z(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0406_),
    .Z(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_14.mux_l1_in_0_.out ),
    .TE_B(_0407_),
    .Z(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0408_),
    .Z(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0409_),
    .Z(\sb_0__0_.mux_right_track_14.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0410_),
    .Z(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0411_),
    .Z(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0412_),
    .Z(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_right_track_2.mux_l1_in_0_.out ),
    .TE_B(_0413_),
    .Z(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0414_),
    .Z(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0415_),
    .Z(\sb_0__0_.mux_right_track_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0416_),
    .Z(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0417_),
    .Z(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0418_),
    .Z(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_top_track_0.mux_l1_in_0_.out ),
    .TE_B(_0419_),
    .Z(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.out ),
    .TE_B(_0420_),
    .Z(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0421_),
    .Z(\sb_0__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0422_),
    .Z(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0423_),
    .Z(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0424_),
    .Z(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__0_.mux_top_track_12.mux_l1_in_0_.out ),
    .TE_B(_0425_),
    .Z(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.out ),
    .TE_B(_0426_),
    .Z(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0427_),
    .Z(\sb_0__0_.mux_top_track_12.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_5.INVTX1_5_.out ),
    .TE_B(_0428_),
    .Z(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0429_),
    .Z(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0430_),
    .Z(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_bottom_track_1.mux_l1_in_0_.out ),
    .TE_B(_0431_),
    .Z(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0432_),
    .Z(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0433_),
    .Z(\sb_0__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_3_.out ),
    .TE_B(_0434_),
    .Z(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0435_),
    .Z(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0436_),
    .Z(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_bottom_track_15.mux_l1_in_0_.out ),
    .TE_B(_0437_),
    .Z(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0438_),
    .Z(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0439_),
    .Z(\sb_0__1_.mux_bottom_track_15.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_4.INVTX1_5_.out ),
    .TE_B(_0440_),
    .Z(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0441_),
    .Z(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0442_),
    .Z(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_bottom_track_3.mux_l1_in_0_.out ),
    .TE_B(_0443_),
    .Z(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0444_),
    .Z(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0445_),
    .Z(\sb_0__1_.mux_bottom_track_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0725_),
    .Z(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0725_),
    .Z(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0725_),
    .Z(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_right_track_0.mux_l1_in_0_.out ),
    .TE_B(_0725_),
    .Z(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_4_.out ),
    .TE_B(_0725_),
    .Z(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0725_),
    .Z(\sb_0__1_.mux_right_track_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0446_),
    .Z(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0447_),
    .Z(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0448_),
    .Z(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_0__1_.mux_right_track_12.mux_l1_in_0_.out ),
    .TE_B(_0449_),
    .Z(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cby_0__1_.mux_right_ipin_3.INVTX1_2_.out ),
    .TE_B(_0450_),
    .Z(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0451_),
    .Z(\sb_0__1_.mux_right_track_12.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.out ),
    .TE_B(_0452_),
    .Z(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0453_),
    .Z(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0454_),
    .Z(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_1.mux_l1_in_0_.out ),
    .TE_B(_0455_),
    .Z(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0456_),
    .Z(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0457_),
    .Z(\sb_1__0_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_1.INVTX1_5_.out ),
    .TE_B(_0458_),
    .Z(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0459_),
    .Z(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0460_),
    .Z(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_13.mux_l1_in_0_.out ),
    .TE_B(_0461_),
    .Z(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0462_),
    .Z(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0463_),
    .Z(\sb_1__0_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.out ),
    .TE_B(_0464_),
    .Z(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0465_),
    .Z(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0466_),
    .Z(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_15.mux_l1_in_0_.out ),
    .TE_B(_0467_),
    .Z(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0468_),
    .Z(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0469_),
    .Z(\sb_1__0_.mux_left_track_15.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_5_.out ),
    .TE_B(_0470_),
    .Z(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0471_),
    .Z(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0472_),
    .Z(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_left_track_3.mux_l1_in_0_.out ),
    .TE_B(_0473_),
    .Z(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0474_),
    .Z(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0475_),
    .Z(\sb_1__0_.mux_left_track_3.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.ble4_0.mux_ble4_out_0.mux_l1_in_0_.out ),
    .TE_B(_0476_),
    .Z(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0477_),
    .Z(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0478_),
    .Z(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_0.mux_l1_in_0_.out ),
    .TE_B(_0479_),
    .Z(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\sb_0__0_.mux_right_track_0.mux_l2_in_0_.out ),
    .TE_B(_0480_),
    .Z(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0481_),
    .Z(\sb_1__0_.mux_top_track_0.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0482_),
    .Z(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0483_),
    .Z(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0484_),
    .Z(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_14.mux_l1_in_0_.out ),
    .TE_B(_0485_),
    .Z(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\sb_0__0_.mux_right_track_12.mux_l2_in_0_.out ),
    .TE_B(_0486_),
    .Z(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0487_),
    .Z(\sb_1__0_.mux_top_track_14.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0488_),
    .Z(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0489_),
    .Z(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0490_),
    .Z(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__0_.mux_top_track_2.mux_l1_in_0_.out ),
    .TE_B(_0491_),
    .Z(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__0_.mux_bottom_ipin_0.INVTX1_4_.out ),
    .TE_B(_0492_),
    .Z(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0493_),
    .Z(\sb_1__0_.mux_top_track_2.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0494_),
    .Z(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0495_),
    .Z(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0496_),
    .Z(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_bottom_track_1.mux_l1_in_0_.out ),
    .TE_B(_0497_),
    .Z(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0498_),
    .Z(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0499_),
    .Z(\sb_1__1_.mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.ebufn  (.A(_0725_),
    .TE_B(_0500_),
    .Z(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0501_),
    .Z(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0502_),
    .Z(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_bottom_track_13.mux_l1_in_0_.out ),
    .TE_B(_0503_),
    .Z(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.ebufn  (.A(\cbx_1__1_.mux_bottom_ipin_1.INVTX1_4_.out ),
    .TE_B(_0504_),
    .Z(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0505_),
    .Z(\sb_1__1_.mux_bottom_track_13.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_0.INVTX1_4_.out ),
    .TE_B(_0506_),
    .Z(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0507_),
    .Z(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0508_),
    .Z(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_left_track_1.mux_l1_in_0_.out ),
    .TE_B(_0509_),
    .Z(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0510_),
    .Z(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0511_),
    .Z(\sb_1__1_.mux_left_track_1.mux_l2_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.ebufn  (.A(\cby_1__1_.mux_left_ipin_5.INVTX1_2_.out ),
    .TE_B(_0512_),
    .Z(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0513_),
    .Z(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0514_),
    .Z(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.TGATE_2_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.ebufn  (.A(\sb_1__1_.mux_left_track_13.mux_l1_in_0_.out ),
    .TE_B(_0515_),
    .Z(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_0_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.ebufn  (.A(_0725_),
    .TE_B(_0516_),
    .Z(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_1_.out ));
 sky130_fd_sc_hd__ebufn_1 \sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.ebufn  (.A(_0725_),
    .TE_B(_0517_),
    .Z(\sb_1__1_.mux_left_track_13.mux_l2_in_0_.TGATE_2_.out ));
endmodule
