VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rram_28
  CLASS BLOCK ;
  FOREIGN rram_28 ;
  ORIGIN 0.330 0.165 ;
  SIZE 23.340 BY 11.525 ;
  PIN Q[2]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 1.985 9.040 2.155 10.770 ;
      LAYER mcon ;
        RECT 1.985 9.605 2.155 9.775 ;
      LAYER met1 ;
        RECT 1.920 9.540 2.520 9.860 ;
      LAYER via ;
        RECT 2.250 9.570 2.510 9.830 ;
      LAYER met2 ;
        RECT 2.240 9.860 2.440 11.360 ;
        RECT 2.240 9.540 2.520 9.860 ;
    END
  END Q[2]
  PIN Q[6]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 5.225 9.040 5.395 10.770 ;
      LAYER mcon ;
        RECT 5.225 9.605 5.395 9.775 ;
      LAYER met1 ;
        RECT 5.160 9.540 5.760 9.860 ;
      LAYER via ;
        RECT 5.490 9.570 5.750 9.830 ;
      LAYER met2 ;
        RECT 5.480 9.860 5.680 11.360 ;
        RECT 5.480 9.540 5.760 9.860 ;
    END
  END Q[6]
  PIN Q[10]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 8.465 9.040 8.635 10.770 ;
      LAYER mcon ;
        RECT 8.465 9.605 8.635 9.775 ;
      LAYER met1 ;
        RECT 8.400 9.540 9.000 9.860 ;
      LAYER via ;
        RECT 8.730 9.570 8.990 9.830 ;
      LAYER met2 ;
        RECT 8.720 9.860 8.920 11.360 ;
        RECT 8.720 9.540 9.000 9.860 ;
    END
  END Q[10]
  PIN Q[18]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 14.945 9.040 15.115 10.770 ;
      LAYER mcon ;
        RECT 14.945 9.605 15.115 9.775 ;
      LAYER met1 ;
        RECT 14.880 9.540 15.480 9.860 ;
      LAYER via ;
        RECT 15.210 9.570 15.470 9.830 ;
      LAYER met2 ;
        RECT 15.200 9.860 15.400 11.360 ;
        RECT 15.200 9.540 15.480 9.860 ;
    END
  END Q[18]
  PIN Q[22]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 18.185 9.040 18.355 10.770 ;
      LAYER mcon ;
        RECT 18.185 9.605 18.355 9.775 ;
      LAYER met1 ;
        RECT 18.120 9.540 18.720 9.860 ;
      LAYER via ;
        RECT 18.450 9.570 18.710 9.830 ;
      LAYER met2 ;
        RECT 18.440 9.860 18.640 11.360 ;
        RECT 18.440 9.540 18.720 9.860 ;
    END
  END Q[22]
  PIN BL[0]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 0.750 7.840 1.230 8.090 ;
      LAYER mcon ;
        RECT 0.900 7.875 1.070 8.045 ;
      LAYER met1 ;
        RECT 0.220 7.790 1.180 8.090 ;
      LAYER via ;
        RECT 0.310 7.810 0.570 8.070 ;
      LAYER met2 ;
        RECT 0.310 7.010 0.570 11.120 ;
        RECT 0.310 0.000 0.570 6.750 ;
    END
  END BL[0]
  PIN BL[4]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 3.990 7.840 4.470 8.090 ;
      LAYER mcon ;
        RECT 4.140 7.875 4.310 8.045 ;
      LAYER met1 ;
        RECT 3.460 7.790 4.420 8.090 ;
      LAYER via ;
        RECT 3.550 7.810 3.810 8.070 ;
      LAYER met2 ;
        RECT 3.550 7.010 3.810 11.120 ;
        RECT 3.550 0.000 3.810 6.750 ;
    END
  END BL[4]
  PIN BL[8]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 7.230 7.840 7.710 8.090 ;
      LAYER mcon ;
        RECT 7.380 7.875 7.550 8.045 ;
      LAYER met1 ;
        RECT 6.700 7.790 7.660 8.090 ;
      LAYER via ;
        RECT 6.790 7.810 7.050 8.070 ;
      LAYER met2 ;
        RECT 6.790 7.010 7.050 11.120 ;
        RECT 6.790 0.000 7.050 6.750 ;
    END
  END BL[8]
  PIN BL[12]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 10.470 7.840 10.950 8.090 ;
      LAYER mcon ;
        RECT 10.620 7.875 10.790 8.045 ;
      LAYER met1 ;
        RECT 9.940 7.790 10.900 8.090 ;
      LAYER via ;
        RECT 10.030 7.810 10.290 8.070 ;
      LAYER met2 ;
        RECT 10.030 7.010 10.290 11.120 ;
        RECT 10.030 0.000 10.290 6.750 ;
    END
  END BL[12]
  PIN BL[16]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 13.710 7.840 14.190 8.090 ;
      LAYER mcon ;
        RECT 13.860 7.875 14.030 8.045 ;
      LAYER met1 ;
        RECT 13.180 7.790 14.140 8.090 ;
      LAYER via ;
        RECT 13.270 7.810 13.530 8.070 ;
      LAYER met2 ;
        RECT 13.270 7.010 13.530 11.120 ;
        RECT 13.270 0.000 13.530 6.750 ;
    END
  END BL[16]
  PIN BL[20]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 16.950 7.840 17.430 8.090 ;
      LAYER mcon ;
        RECT 17.100 7.875 17.270 8.045 ;
      LAYER met1 ;
        RECT 16.420 7.790 17.380 8.090 ;
      LAYER via ;
        RECT 16.510 7.810 16.770 8.070 ;
      LAYER met2 ;
        RECT 16.510 7.010 16.770 11.120 ;
        RECT 16.510 0.000 16.770 6.750 ;
    END
  END BL[20]
  PIN BL[24]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 20.190 7.840 20.670 8.090 ;
      LAYER mcon ;
        RECT 20.340 7.875 20.510 8.045 ;
      LAYER met1 ;
        RECT 19.660 7.790 20.620 8.090 ;
      LAYER via ;
        RECT 19.750 7.810 20.010 8.070 ;
      LAYER met2 ;
        RECT 19.750 7.010 20.010 11.120 ;
        RECT 19.750 0.000 20.010 6.750 ;
    END
  END BL[24]
  PIN BL[1]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 0.530 3.210 1.010 3.460 ;
      LAYER mcon ;
        RECT 0.690 3.255 0.860 3.425 ;
      LAYER met1 ;
        RECT 0.580 3.210 1.540 3.510 ;
      LAYER via ;
        RECT 1.190 3.230 1.450 3.490 ;
      LAYER met2 ;
        RECT 1.190 4.510 1.450 11.120 ;
        RECT 1.190 0.000 1.450 4.250 ;
    END
  END BL[1]
  PIN BL[5]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 3.770 3.210 4.250 3.460 ;
      LAYER mcon ;
        RECT 3.930 3.255 4.100 3.425 ;
      LAYER met1 ;
        RECT 3.820 3.210 4.780 3.510 ;
      LAYER via ;
        RECT 4.430 3.230 4.690 3.490 ;
      LAYER met2 ;
        RECT 4.430 4.510 4.690 11.120 ;
        RECT 4.430 0.000 4.690 4.250 ;
    END
  END BL[5]
  PIN BL[9]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 7.010 3.210 7.490 3.460 ;
      LAYER mcon ;
        RECT 7.170 3.255 7.340 3.425 ;
      LAYER met1 ;
        RECT 7.060 3.210 8.020 3.510 ;
      LAYER via ;
        RECT 7.670 3.230 7.930 3.490 ;
      LAYER met2 ;
        RECT 7.670 4.510 7.930 11.120 ;
        RECT 7.670 0.000 7.930 4.250 ;
    END
  END BL[9]
  PIN BL[13]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 10.250 3.210 10.730 3.460 ;
      LAYER mcon ;
        RECT 10.410 3.255 10.580 3.425 ;
      LAYER met1 ;
        RECT 10.300 3.210 11.260 3.510 ;
      LAYER via ;
        RECT 10.910 3.230 11.170 3.490 ;
      LAYER met2 ;
        RECT 10.910 4.510 11.170 11.120 ;
        RECT 10.910 0.000 11.170 4.250 ;
    END
  END BL[13]
  PIN BL[17]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 13.490 3.210 13.970 3.460 ;
      LAYER mcon ;
        RECT 13.650 3.255 13.820 3.425 ;
      LAYER met1 ;
        RECT 13.540 3.210 14.500 3.510 ;
      LAYER via ;
        RECT 14.150 3.230 14.410 3.490 ;
      LAYER met2 ;
        RECT 14.150 4.510 14.410 11.120 ;
        RECT 14.150 0.000 14.410 4.250 ;
    END
  END BL[17]
  PIN BL[21]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 16.730 3.210 17.210 3.460 ;
      LAYER mcon ;
        RECT 16.890 3.255 17.060 3.425 ;
      LAYER met1 ;
        RECT 16.780 3.210 17.740 3.510 ;
      LAYER via ;
        RECT 17.390 3.230 17.650 3.490 ;
      LAYER met2 ;
        RECT 17.390 4.510 17.650 11.120 ;
        RECT 17.390 0.000 17.650 4.250 ;
    END
  END BL[21]
  PIN BL[25]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 19.970 3.210 20.450 3.460 ;
      LAYER mcon ;
        RECT 20.130 3.255 20.300 3.425 ;
      LAYER met1 ;
        RECT 20.020 3.210 20.980 3.510 ;
      LAYER via ;
        RECT 20.630 3.230 20.890 3.490 ;
      LAYER met2 ;
        RECT 20.630 4.510 20.890 11.120 ;
        RECT 20.630 0.000 20.890 4.250 ;
    END
  END BL[25]
  PIN BL[2]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 2.230 7.840 2.710 8.090 ;
      LAYER mcon ;
        RECT 2.380 7.875 2.550 8.045 ;
      LAYER met1 ;
        RECT 1.700 7.790 2.660 8.090 ;
      LAYER via ;
        RECT 1.790 7.810 2.050 8.070 ;
      LAYER met2 ;
        RECT 1.790 7.010 2.050 11.120 ;
        RECT 1.790 0.000 2.050 6.750 ;
    END
  END BL[2]
  PIN BL[6]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 5.470 7.840 5.950 8.090 ;
      LAYER mcon ;
        RECT 5.620 7.875 5.790 8.045 ;
      LAYER met1 ;
        RECT 4.940 7.790 5.900 8.090 ;
      LAYER via ;
        RECT 5.030 7.810 5.290 8.070 ;
      LAYER met2 ;
        RECT 5.030 7.010 5.290 11.120 ;
        RECT 5.030 0.000 5.290 6.750 ;
    END
  END BL[6]
  PIN BL[10]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 8.710 7.840 9.190 8.090 ;
      LAYER mcon ;
        RECT 8.860 7.875 9.030 8.045 ;
      LAYER met1 ;
        RECT 8.180 7.790 9.140 8.090 ;
      LAYER via ;
        RECT 8.270 7.810 8.530 8.070 ;
      LAYER met2 ;
        RECT 8.270 7.010 8.530 11.120 ;
        RECT 8.270 0.000 8.530 6.750 ;
    END
  END BL[10]
  PIN BL[14]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 11.950 7.840 12.430 8.090 ;
      LAYER mcon ;
        RECT 12.100 7.875 12.270 8.045 ;
      LAYER met1 ;
        RECT 11.420 7.790 12.380 8.090 ;
      LAYER via ;
        RECT 11.510 7.810 11.770 8.070 ;
      LAYER met2 ;
        RECT 11.510 7.010 11.770 11.120 ;
        RECT 11.510 0.000 11.770 6.750 ;
    END
  END BL[14]
  PIN BL[18]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 15.190 7.840 15.670 8.090 ;
      LAYER mcon ;
        RECT 15.340 7.875 15.510 8.045 ;
      LAYER met1 ;
        RECT 14.660 7.790 15.620 8.090 ;
      LAYER via ;
        RECT 14.750 7.810 15.010 8.070 ;
      LAYER met2 ;
        RECT 14.750 7.010 15.010 11.120 ;
        RECT 14.750 0.000 15.010 6.750 ;
    END
  END BL[18]
  PIN BL[22]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 18.430 7.840 18.910 8.090 ;
      LAYER mcon ;
        RECT 18.580 7.875 18.750 8.045 ;
      LAYER met1 ;
        RECT 17.900 7.790 18.860 8.090 ;
      LAYER via ;
        RECT 17.990 7.810 18.250 8.070 ;
      LAYER met2 ;
        RECT 17.990 7.010 18.250 11.120 ;
        RECT 17.990 0.000 18.250 6.750 ;
    END
  END BL[22]
  PIN BL[26]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 21.670 7.840 22.150 8.090 ;
      LAYER mcon ;
        RECT 21.820 7.875 21.990 8.045 ;
      LAYER met1 ;
        RECT 21.140 7.790 22.100 8.090 ;
      LAYER via ;
        RECT 21.230 7.810 21.490 8.070 ;
      LAYER met2 ;
        RECT 21.230 7.010 21.490 11.120 ;
        RECT 21.230 0.000 21.490 6.750 ;
    END
  END BL[26]
  PIN BL[3]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 2.010 3.210 2.490 3.460 ;
      LAYER mcon ;
        RECT 2.170 3.255 2.340 3.425 ;
      LAYER met1 ;
        RECT 2.060 3.210 3.020 3.510 ;
      LAYER via ;
        RECT 2.670 3.230 2.930 3.490 ;
      LAYER met2 ;
        RECT 2.670 4.510 2.930 11.120 ;
        RECT 2.670 0.000 2.930 4.250 ;
    END
  END BL[3]
  PIN BL[7]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 5.250 3.210 5.730 3.460 ;
      LAYER mcon ;
        RECT 5.410 3.255 5.580 3.425 ;
      LAYER met1 ;
        RECT 5.300 3.210 6.260 3.510 ;
      LAYER via ;
        RECT 5.910 3.230 6.170 3.490 ;
      LAYER met2 ;
        RECT 5.910 4.510 6.170 11.120 ;
        RECT 5.910 0.000 6.170 4.250 ;
    END
  END BL[7]
  PIN BL[11]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 8.490 3.210 8.970 3.460 ;
      LAYER mcon ;
        RECT 8.650 3.255 8.820 3.425 ;
      LAYER met1 ;
        RECT 8.540 3.210 9.500 3.510 ;
      LAYER via ;
        RECT 9.150 3.230 9.410 3.490 ;
      LAYER met2 ;
        RECT 9.150 4.510 9.410 11.120 ;
        RECT 9.150 0.000 9.410 4.250 ;
    END
  END BL[11]
  PIN BL[15]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 11.730 3.210 12.210 3.460 ;
      LAYER mcon ;
        RECT 11.890 3.255 12.060 3.425 ;
      LAYER met1 ;
        RECT 11.780 3.210 12.740 3.510 ;
      LAYER via ;
        RECT 12.390 3.230 12.650 3.490 ;
      LAYER met2 ;
        RECT 12.390 4.510 12.650 11.120 ;
        RECT 12.390 0.000 12.650 4.250 ;
    END
  END BL[15]
  PIN BL[19]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 14.970 3.210 15.450 3.460 ;
      LAYER mcon ;
        RECT 15.130 3.255 15.300 3.425 ;
      LAYER met1 ;
        RECT 15.020 3.210 15.980 3.510 ;
      LAYER via ;
        RECT 15.630 3.230 15.890 3.490 ;
      LAYER met2 ;
        RECT 15.630 4.510 15.890 11.120 ;
        RECT 15.630 0.000 15.890 4.250 ;
    END
  END BL[19]
  PIN BL[23]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 18.210 3.210 18.690 3.460 ;
      LAYER mcon ;
        RECT 18.370 3.255 18.540 3.425 ;
      LAYER met1 ;
        RECT 18.260 3.210 19.220 3.510 ;
      LAYER via ;
        RECT 18.870 3.230 19.130 3.490 ;
      LAYER met2 ;
        RECT 18.870 4.510 19.130 11.120 ;
        RECT 18.870 0.000 19.130 4.250 ;
    END
  END BL[23]
  PIN BL[27]
    ANTENNAGATEAREA 0.750000 ;
    PORT
      LAYER li1 ;
        RECT 21.450 3.210 21.930 3.460 ;
      LAYER mcon ;
        RECT 21.610 3.255 21.780 3.425 ;
      LAYER met1 ;
        RECT 21.500 3.210 22.460 3.510 ;
      LAYER via ;
        RECT 22.110 3.230 22.370 3.490 ;
      LAYER met2 ;
        RECT 22.110 4.510 22.370 11.120 ;
        RECT 22.110 0.000 22.370 4.250 ;
    END
  END BL[27]
  PIN Q[0]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 0.385 9.040 0.555 10.790 ;
      LAYER mcon ;
        RECT 0.385 9.605 0.555 9.775 ;
      LAYER met1 ;
        RECT 0.320 9.540 1.040 9.880 ;
      LAYER via ;
        RECT 0.770 9.570 1.030 9.830 ;
      LAYER met2 ;
        RECT 0.750 9.880 0.950 11.360 ;
        RECT 0.750 9.540 1.040 9.880 ;
    END
  END Q[0]
  PIN Q[4]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 3.625 9.040 3.795 10.790 ;
      LAYER mcon ;
        RECT 3.625 9.605 3.795 9.775 ;
      LAYER met1 ;
        RECT 3.560 9.540 4.280 9.880 ;
      LAYER via ;
        RECT 4.010 9.570 4.270 9.830 ;
      LAYER met2 ;
        RECT 3.990 9.880 4.190 11.360 ;
        RECT 3.990 9.540 4.280 9.880 ;
    END
  END Q[4]
  PIN Q[8]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 6.865 9.040 7.035 10.790 ;
      LAYER mcon ;
        RECT 6.865 9.605 7.035 9.775 ;
      LAYER met1 ;
        RECT 6.800 9.540 7.520 9.880 ;
      LAYER via ;
        RECT 7.250 9.570 7.510 9.830 ;
      LAYER met2 ;
        RECT 7.230 9.880 7.430 11.360 ;
        RECT 7.230 9.540 7.520 9.880 ;
    END
  END Q[8]
  PIN Q[12]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 10.105 9.040 10.275 10.790 ;
      LAYER mcon ;
        RECT 10.105 9.605 10.275 9.775 ;
      LAYER met1 ;
        RECT 10.040 9.540 10.760 9.880 ;
      LAYER via ;
        RECT 10.490 9.570 10.750 9.830 ;
      LAYER met2 ;
        RECT 10.470 9.880 10.670 11.360 ;
        RECT 10.470 9.540 10.760 9.880 ;
    END
  END Q[12]
  PIN Q[16]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 13.345 9.040 13.515 10.790 ;
      LAYER mcon ;
        RECT 13.345 9.605 13.515 9.775 ;
      LAYER met1 ;
        RECT 13.280 9.540 14.000 9.880 ;
      LAYER via ;
        RECT 13.730 9.570 13.990 9.830 ;
      LAYER met2 ;
        RECT 13.710 9.880 13.910 11.360 ;
        RECT 13.710 9.540 14.000 9.880 ;
    END
  END Q[16]
  PIN Q[20]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 16.585 9.040 16.755 10.790 ;
      LAYER mcon ;
        RECT 16.585 9.605 16.755 9.775 ;
      LAYER met1 ;
        RECT 16.520 9.540 17.240 9.880 ;
      LAYER via ;
        RECT 16.970 9.570 17.230 9.830 ;
      LAYER met2 ;
        RECT 16.950 9.880 17.150 11.360 ;
        RECT 16.950 9.540 17.240 9.880 ;
    END
  END Q[20]
  PIN Q[24]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 19.825 9.040 19.995 10.790 ;
      LAYER mcon ;
        RECT 19.825 9.605 19.995 9.775 ;
      LAYER met1 ;
        RECT 19.760 9.540 20.480 9.880 ;
      LAYER via ;
        RECT 20.210 9.570 20.470 9.830 ;
      LAYER met2 ;
        RECT 20.190 9.880 20.390 11.360 ;
        RECT 20.190 9.540 20.480 9.880 ;
    END
  END Q[24]
  PIN Q[14]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 11.705 9.040 11.875 10.770 ;
      LAYER mcon ;
        RECT 11.705 9.605 11.875 9.775 ;
      LAYER met1 ;
        RECT 11.640 9.540 12.240 9.860 ;
      LAYER via ;
        RECT 11.970 9.570 12.230 9.830 ;
      LAYER met2 ;
        RECT 11.960 9.860 12.160 11.360 ;
        RECT 11.960 9.540 12.240 9.860 ;
    END
  END Q[14]
  PIN Q[26]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 21.425 9.040 21.595 10.770 ;
      LAYER mcon ;
        RECT 21.425 9.605 21.595 9.775 ;
      LAYER met1 ;
        RECT 21.360 9.540 21.960 9.860 ;
      LAYER via ;
        RECT 21.690 9.570 21.950 9.830 ;
      LAYER met2 ;
        RECT 21.680 9.860 21.880 11.360 ;
        RECT 21.680 9.540 21.960 9.860 ;
    END
  END Q[26]
  PIN Q[1]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 1.085 0.590 1.255 2.320 ;
      LAYER mcon ;
        RECT 1.085 1.585 1.255 1.755 ;
      LAYER met1 ;
        RECT 0.720 1.500 1.320 1.820 ;
      LAYER via ;
        RECT 0.730 1.530 0.990 1.790 ;
      LAYER met2 ;
        RECT 0.720 1.500 1.000 1.820 ;
        RECT 0.800 0.000 1.000 1.500 ;
    END
  END Q[1]
  PIN Q[5]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 4.325 0.590 4.495 2.320 ;
      LAYER mcon ;
        RECT 4.325 1.585 4.495 1.755 ;
      LAYER met1 ;
        RECT 3.960 1.500 4.560 1.820 ;
      LAYER via ;
        RECT 3.970 1.530 4.230 1.790 ;
      LAYER met2 ;
        RECT 3.960 1.500 4.240 1.820 ;
        RECT 4.040 0.000 4.240 1.500 ;
    END
  END Q[5]
  PIN Q[13]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 10.805 0.590 10.975 2.320 ;
      LAYER mcon ;
        RECT 10.805 1.585 10.975 1.755 ;
      LAYER met1 ;
        RECT 10.440 1.500 11.040 1.820 ;
      LAYER via ;
        RECT 10.450 1.530 10.710 1.790 ;
      LAYER met2 ;
        RECT 10.440 1.500 10.720 1.820 ;
        RECT 10.520 0.000 10.720 1.500 ;
    END
  END Q[13]
  PIN Q[17]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 14.045 0.590 14.215 2.320 ;
      LAYER mcon ;
        RECT 14.045 1.585 14.215 1.755 ;
      LAYER met1 ;
        RECT 13.680 1.500 14.280 1.820 ;
      LAYER via ;
        RECT 13.690 1.530 13.950 1.790 ;
      LAYER met2 ;
        RECT 13.680 1.500 13.960 1.820 ;
        RECT 13.760 0.000 13.960 1.500 ;
    END
  END Q[17]
  PIN Q[21]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 17.285 0.590 17.455 2.320 ;
      LAYER mcon ;
        RECT 17.285 1.585 17.455 1.755 ;
      LAYER met1 ;
        RECT 16.920 1.500 17.520 1.820 ;
      LAYER via ;
        RECT 16.930 1.530 17.190 1.790 ;
      LAYER met2 ;
        RECT 16.920 1.500 17.200 1.820 ;
        RECT 17.000 0.000 17.200 1.500 ;
    END
  END Q[21]
  PIN Q[25]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 20.525 0.590 20.695 2.320 ;
      LAYER mcon ;
        RECT 20.525 1.585 20.695 1.755 ;
      LAYER met1 ;
        RECT 20.160 1.500 20.760 1.820 ;
      LAYER via ;
        RECT 20.170 1.530 20.430 1.790 ;
      LAYER met2 ;
        RECT 20.160 1.500 20.440 1.820 ;
        RECT 20.240 0.000 20.440 1.500 ;
    END
  END Q[25]
  PIN Q[9]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 7.565 0.590 7.735 2.320 ;
      LAYER mcon ;
        RECT 7.565 1.585 7.735 1.755 ;
      LAYER met1 ;
        RECT 7.200 1.500 7.800 1.820 ;
      LAYER via ;
        RECT 7.210 1.530 7.470 1.790 ;
      LAYER met2 ;
        RECT 7.200 1.500 7.480 1.820 ;
        RECT 7.280 0.000 7.480 1.500 ;
    END
  END Q[9]
  PIN Q[3]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 2.685 0.570 2.855 2.320 ;
      LAYER mcon ;
        RECT 2.685 1.585 2.855 1.755 ;
      LAYER met1 ;
        RECT 2.200 1.480 2.920 1.820 ;
      LAYER via ;
        RECT 2.210 1.530 2.470 1.790 ;
      LAYER met2 ;
        RECT 2.200 1.480 2.490 1.820 ;
        RECT 2.290 0.000 2.490 1.480 ;
    END
  END Q[3]
  PIN Q[7]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 5.925 0.570 6.095 2.320 ;
      LAYER mcon ;
        RECT 5.925 1.585 6.095 1.755 ;
      LAYER met1 ;
        RECT 5.440 1.480 6.160 1.820 ;
      LAYER via ;
        RECT 5.450 1.530 5.710 1.790 ;
      LAYER met2 ;
        RECT 5.440 1.480 5.730 1.820 ;
        RECT 5.530 0.000 5.730 1.480 ;
    END
  END Q[7]
  PIN Q[15]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 12.405 0.570 12.575 2.320 ;
      LAYER mcon ;
        RECT 12.405 1.585 12.575 1.755 ;
      LAYER met1 ;
        RECT 11.920 1.480 12.640 1.820 ;
      LAYER via ;
        RECT 11.930 1.530 12.190 1.790 ;
      LAYER met2 ;
        RECT 11.920 1.480 12.210 1.820 ;
        RECT 12.010 0.000 12.210 1.480 ;
    END
  END Q[15]
  PIN Q[19]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 15.645 0.570 15.815 2.320 ;
      LAYER mcon ;
        RECT 15.645 1.585 15.815 1.755 ;
      LAYER met1 ;
        RECT 15.160 1.480 15.880 1.820 ;
      LAYER via ;
        RECT 15.170 1.530 15.430 1.790 ;
      LAYER met2 ;
        RECT 15.160 1.480 15.450 1.820 ;
        RECT 15.250 0.000 15.450 1.480 ;
    END
  END Q[19]
  PIN Q[23]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 18.885 0.570 19.055 2.320 ;
      LAYER mcon ;
        RECT 18.885 1.585 19.055 1.755 ;
      LAYER met1 ;
        RECT 18.400 1.480 19.120 1.820 ;
      LAYER via ;
        RECT 18.410 1.530 18.670 1.790 ;
      LAYER met2 ;
        RECT 18.400 1.480 18.690 1.820 ;
        RECT 18.490 0.000 18.690 1.480 ;
    END
  END Q[23]
  PIN Q[27]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 22.125 0.570 22.295 2.320 ;
      LAYER mcon ;
        RECT 22.125 1.585 22.295 1.755 ;
      LAYER met1 ;
        RECT 21.640 1.480 22.360 1.820 ;
      LAYER via ;
        RECT 21.650 1.530 21.910 1.790 ;
      LAYER met2 ;
        RECT 21.640 1.480 21.930 1.820 ;
        RECT 21.730 0.000 21.930 1.480 ;
    END
  END Q[27]
  PIN Q[11]
    ANTENNADIFFAREA 0.365400 ;
    PORT
      LAYER li1 ;
        RECT 9.165 0.570 9.335 2.320 ;
      LAYER mcon ;
        RECT 9.165 1.585 9.335 1.755 ;
      LAYER met1 ;
        RECT 8.680 1.480 9.400 1.820 ;
      LAYER via ;
        RECT 8.690 1.530 8.950 1.790 ;
      LAYER met2 ;
        RECT 8.680 1.480 8.970 1.820 ;
        RECT 8.770 0.000 8.970 1.480 ;
    END
  END Q[11]
  OBS
      LAYER nwell ;
        RECT 0.000 9.800 22.680 11.260 ;
      LAYER pwell ;
        RECT 1.265 9.590 1.695 9.775 ;
        RECT 4.505 9.590 4.935 9.775 ;
        RECT 7.745 9.590 8.175 9.775 ;
        RECT 10.985 9.590 11.415 9.775 ;
        RECT 14.225 9.590 14.655 9.775 ;
        RECT 17.465 9.590 17.895 9.775 ;
        RECT 20.705 9.590 21.135 9.775 ;
        RECT 0.195 8.910 2.785 9.590 ;
        RECT 3.435 8.910 6.025 9.590 ;
        RECT 6.675 8.910 9.265 9.590 ;
        RECT 9.915 8.910 12.505 9.590 ;
        RECT 13.155 8.910 15.745 9.590 ;
        RECT 16.395 8.910 18.985 9.590 ;
        RECT 19.635 8.910 22.225 9.590 ;
        RECT 0.965 8.715 1.135 8.910 ;
        RECT 4.205 8.715 4.375 8.910 ;
        RECT 7.445 8.715 7.615 8.910 ;
        RECT 10.685 8.715 10.855 8.910 ;
        RECT 13.925 8.715 14.095 8.910 ;
        RECT 17.165 8.715 17.335 8.910 ;
        RECT 20.405 8.715 20.575 8.910 ;
      LAYER nwell ;
        RECT -0.330 3.320 23.010 8.120 ;
      LAYER pwell ;
        RECT 2.105 2.450 2.275 2.645 ;
        RECT 5.345 2.450 5.515 2.645 ;
        RECT 8.585 2.450 8.755 2.645 ;
        RECT 11.825 2.450 11.995 2.645 ;
        RECT 15.065 2.450 15.235 2.645 ;
        RECT 18.305 2.450 18.475 2.645 ;
        RECT 21.545 2.450 21.715 2.645 ;
        RECT 0.455 1.770 3.045 2.450 ;
        RECT 3.695 1.770 6.285 2.450 ;
        RECT 6.935 1.770 9.525 2.450 ;
        RECT 10.175 1.770 12.765 2.450 ;
        RECT 13.415 1.770 16.005 2.450 ;
        RECT 16.655 1.770 19.245 2.450 ;
        RECT 19.895 1.770 22.485 2.450 ;
        RECT 1.545 1.585 1.975 1.770 ;
        RECT 4.785 1.585 5.215 1.770 ;
        RECT 8.025 1.585 8.455 1.770 ;
        RECT 11.265 1.585 11.695 1.770 ;
        RECT 14.505 1.585 14.935 1.770 ;
        RECT 17.745 1.585 18.175 1.770 ;
        RECT 20.985 1.585 21.415 1.770 ;
      LAYER nwell ;
        RECT 0.000 0.100 22.680 1.560 ;
      LAYER li1 ;
        RECT 0.000 11.035 3.000 11.205 ;
        RECT 3.240 11.035 6.240 11.205 ;
        RECT 6.480 11.035 9.480 11.205 ;
        RECT 9.720 11.035 12.720 11.205 ;
        RECT 12.960 11.035 15.960 11.205 ;
        RECT 16.200 11.035 19.200 11.205 ;
        RECT 19.440 11.035 22.440 11.205 ;
        RECT 0.825 9.990 0.995 11.035 ;
        RECT 2.425 9.990 2.595 11.035 ;
        RECT 4.065 9.990 4.235 11.035 ;
        RECT 5.665 9.990 5.835 11.035 ;
        RECT 7.305 9.990 7.475 11.035 ;
        RECT 8.905 9.990 9.075 11.035 ;
        RECT 10.545 9.990 10.715 11.035 ;
        RECT 12.145 9.990 12.315 11.035 ;
        RECT 13.785 9.990 13.955 11.035 ;
        RECT 15.385 9.990 15.555 11.035 ;
        RECT 17.025 9.990 17.195 11.035 ;
        RECT 18.625 9.990 18.795 11.035 ;
        RECT 20.265 9.990 20.435 11.035 ;
        RECT 21.865 9.990 22.035 11.035 ;
        RECT 0.825 8.885 0.995 9.460 ;
        RECT 1.335 8.885 1.625 9.610 ;
        RECT 2.425 8.885 2.595 9.460 ;
        RECT 4.065 8.885 4.235 9.460 ;
        RECT 4.575 8.885 4.865 9.610 ;
        RECT 5.665 8.885 5.835 9.460 ;
        RECT 7.305 8.885 7.475 9.460 ;
        RECT 7.815 8.885 8.105 9.610 ;
        RECT 8.905 8.885 9.075 9.460 ;
        RECT 10.545 8.885 10.715 9.460 ;
        RECT 11.055 8.885 11.345 9.610 ;
        RECT 12.145 8.885 12.315 9.460 ;
        RECT 13.785 8.885 13.955 9.460 ;
        RECT 14.295 8.885 14.585 9.610 ;
        RECT 15.385 8.885 15.555 9.460 ;
        RECT 17.025 8.885 17.195 9.460 ;
        RECT 17.535 8.885 17.825 9.610 ;
        RECT 18.625 8.885 18.795 9.460 ;
        RECT 20.265 8.885 20.435 9.460 ;
        RECT 20.775 8.885 21.065 9.610 ;
        RECT 21.865 8.885 22.035 9.460 ;
        RECT 0.280 8.620 0.650 8.800 ;
        RECT 0.820 8.715 1.710 8.885 ;
        RECT 1.880 8.620 2.250 8.800 ;
        RECT 2.420 8.715 3.000 8.885 ;
        RECT 3.520 8.620 3.890 8.800 ;
        RECT 4.060 8.715 4.950 8.885 ;
        RECT 5.120 8.620 5.490 8.800 ;
        RECT 5.660 8.715 6.240 8.885 ;
        RECT 6.760 8.620 7.130 8.800 ;
        RECT 7.300 8.715 8.190 8.885 ;
        RECT 8.360 8.620 8.730 8.800 ;
        RECT 8.900 8.715 9.480 8.885 ;
        RECT 10.000 8.620 10.370 8.800 ;
        RECT 10.540 8.715 11.430 8.885 ;
        RECT 11.600 8.620 11.970 8.800 ;
        RECT 12.140 8.715 12.720 8.885 ;
        RECT 13.240 8.620 13.610 8.800 ;
        RECT 13.780 8.715 14.670 8.885 ;
        RECT 14.840 8.620 15.210 8.800 ;
        RECT 15.380 8.715 15.960 8.885 ;
        RECT 16.480 8.620 16.850 8.800 ;
        RECT 17.020 8.715 17.910 8.885 ;
        RECT 18.080 8.620 18.450 8.800 ;
        RECT 18.620 8.715 19.200 8.885 ;
        RECT 19.720 8.620 20.090 8.800 ;
        RECT 20.260 8.715 21.150 8.885 ;
        RECT 21.320 8.620 21.690 8.800 ;
        RECT 21.860 8.715 22.440 8.885 ;
        RECT 0.400 6.120 0.570 8.620 ;
        RECT 1.190 5.940 1.360 7.370 ;
        RECT 1.880 6.120 2.050 8.620 ;
        RECT 2.670 5.940 2.840 7.660 ;
        RECT 3.640 6.120 3.810 8.620 ;
        RECT 4.430 5.940 4.600 7.370 ;
        RECT 5.120 6.120 5.290 8.620 ;
        RECT 5.910 5.940 6.080 7.660 ;
        RECT 6.880 6.120 7.050 8.620 ;
        RECT 7.670 5.940 7.840 7.370 ;
        RECT 8.360 6.120 8.530 8.620 ;
        RECT 9.150 5.940 9.320 7.660 ;
        RECT 10.120 6.120 10.290 8.620 ;
        RECT 10.910 5.940 11.080 7.370 ;
        RECT 11.600 6.120 11.770 8.620 ;
        RECT 12.390 5.940 12.560 7.660 ;
        RECT 13.360 6.120 13.530 8.620 ;
        RECT 14.150 5.940 14.320 7.370 ;
        RECT 14.840 6.120 15.010 8.620 ;
        RECT 15.630 5.940 15.800 7.660 ;
        RECT 16.600 6.120 16.770 8.620 ;
        RECT 17.390 5.940 17.560 7.370 ;
        RECT 18.080 6.120 18.250 8.620 ;
        RECT 18.870 5.940 19.040 7.660 ;
        RECT 19.840 6.120 20.010 8.620 ;
        RECT 20.630 5.940 20.800 7.370 ;
        RECT 21.320 6.120 21.490 8.620 ;
        RECT 22.110 5.940 22.280 7.660 ;
        RECT 0.000 5.360 22.680 5.940 ;
        RECT 0.400 3.740 0.570 5.360 ;
        RECT 1.190 2.740 1.360 5.180 ;
        RECT 1.880 3.750 2.050 5.360 ;
        RECT 2.670 2.740 2.840 5.180 ;
        RECT 3.640 3.740 3.810 5.360 ;
        RECT 4.430 2.740 4.600 5.180 ;
        RECT 5.120 3.750 5.290 5.360 ;
        RECT 5.910 2.740 6.080 5.180 ;
        RECT 6.880 3.740 7.050 5.360 ;
        RECT 7.670 2.740 7.840 5.180 ;
        RECT 8.360 3.750 8.530 5.360 ;
        RECT 9.150 2.740 9.320 5.180 ;
        RECT 10.120 3.740 10.290 5.360 ;
        RECT 10.910 2.740 11.080 5.180 ;
        RECT 11.600 3.750 11.770 5.360 ;
        RECT 12.390 2.740 12.560 5.180 ;
        RECT 13.360 3.740 13.530 5.360 ;
        RECT 14.150 2.740 14.320 5.180 ;
        RECT 14.840 3.750 15.010 5.360 ;
        RECT 15.630 2.740 15.800 5.180 ;
        RECT 16.600 3.740 16.770 5.360 ;
        RECT 17.390 2.740 17.560 5.180 ;
        RECT 18.080 3.750 18.250 5.360 ;
        RECT 18.870 2.740 19.040 5.180 ;
        RECT 19.840 3.740 20.010 5.360 ;
        RECT 20.630 2.740 20.800 5.180 ;
        RECT 21.320 3.750 21.490 5.360 ;
        RECT 22.110 2.740 22.280 5.180 ;
        RECT 0.240 2.475 0.820 2.645 ;
        RECT 0.990 2.560 1.360 2.740 ;
        RECT 1.530 2.475 2.420 2.645 ;
        RECT 2.590 2.560 2.960 2.740 ;
        RECT 3.480 2.475 4.060 2.645 ;
        RECT 4.230 2.560 4.600 2.740 ;
        RECT 4.770 2.475 5.660 2.645 ;
        RECT 5.830 2.560 6.200 2.740 ;
        RECT 6.720 2.475 7.300 2.645 ;
        RECT 7.470 2.560 7.840 2.740 ;
        RECT 8.010 2.475 8.900 2.645 ;
        RECT 9.070 2.560 9.440 2.740 ;
        RECT 9.960 2.475 10.540 2.645 ;
        RECT 10.710 2.560 11.080 2.740 ;
        RECT 11.250 2.475 12.140 2.645 ;
        RECT 12.310 2.560 12.680 2.740 ;
        RECT 13.200 2.475 13.780 2.645 ;
        RECT 13.950 2.560 14.320 2.740 ;
        RECT 14.490 2.475 15.380 2.645 ;
        RECT 15.550 2.560 15.920 2.740 ;
        RECT 16.440 2.475 17.020 2.645 ;
        RECT 17.190 2.560 17.560 2.740 ;
        RECT 17.730 2.475 18.620 2.645 ;
        RECT 18.790 2.560 19.160 2.740 ;
        RECT 19.680 2.475 20.260 2.645 ;
        RECT 20.430 2.560 20.800 2.740 ;
        RECT 20.970 2.475 21.860 2.645 ;
        RECT 22.030 2.560 22.400 2.740 ;
        RECT 0.645 1.900 0.815 2.475 ;
        RECT 1.615 1.750 1.905 2.475 ;
        RECT 2.245 1.900 2.415 2.475 ;
        RECT 3.885 1.900 4.055 2.475 ;
        RECT 4.855 1.750 5.145 2.475 ;
        RECT 5.485 1.900 5.655 2.475 ;
        RECT 7.125 1.900 7.295 2.475 ;
        RECT 8.095 1.750 8.385 2.475 ;
        RECT 8.725 1.900 8.895 2.475 ;
        RECT 10.365 1.900 10.535 2.475 ;
        RECT 11.335 1.750 11.625 2.475 ;
        RECT 11.965 1.900 12.135 2.475 ;
        RECT 13.605 1.900 13.775 2.475 ;
        RECT 14.575 1.750 14.865 2.475 ;
        RECT 15.205 1.900 15.375 2.475 ;
        RECT 16.845 1.900 17.015 2.475 ;
        RECT 17.815 1.750 18.105 2.475 ;
        RECT 18.445 1.900 18.615 2.475 ;
        RECT 20.085 1.900 20.255 2.475 ;
        RECT 21.055 1.750 21.345 2.475 ;
        RECT 21.685 1.900 21.855 2.475 ;
        RECT 0.645 0.325 0.815 1.370 ;
        RECT 2.245 0.325 2.415 1.370 ;
        RECT 3.885 0.325 4.055 1.370 ;
        RECT 5.485 0.325 5.655 1.370 ;
        RECT 7.125 0.325 7.295 1.370 ;
        RECT 8.725 0.325 8.895 1.370 ;
        RECT 10.365 0.325 10.535 1.370 ;
        RECT 11.965 0.325 12.135 1.370 ;
        RECT 13.605 0.325 13.775 1.370 ;
        RECT 15.205 0.325 15.375 1.370 ;
        RECT 16.845 0.325 17.015 1.370 ;
        RECT 18.445 0.325 18.615 1.370 ;
        RECT 20.085 0.325 20.255 1.370 ;
        RECT 21.685 0.325 21.855 1.370 ;
        RECT 0.240 0.155 3.240 0.325 ;
        RECT 3.480 0.155 6.480 0.325 ;
        RECT 6.720 0.155 9.720 0.325 ;
        RECT 9.960 0.155 12.960 0.325 ;
        RECT 13.200 0.155 16.200 0.325 ;
        RECT 16.440 0.155 19.440 0.325 ;
        RECT 19.680 0.155 22.680 0.325 ;
      LAYER mcon ;
        RECT 0.145 11.035 0.315 11.205 ;
        RECT 0.605 11.035 0.775 11.205 ;
        RECT 1.065 11.035 1.235 11.205 ;
        RECT 1.745 11.035 1.915 11.205 ;
        RECT 2.205 11.035 2.375 11.205 ;
        RECT 2.665 11.035 2.835 11.205 ;
        RECT 3.385 11.035 3.555 11.205 ;
        RECT 3.845 11.035 4.015 11.205 ;
        RECT 4.305 11.035 4.475 11.205 ;
        RECT 4.985 11.035 5.155 11.205 ;
        RECT 5.445 11.035 5.615 11.205 ;
        RECT 5.905 11.035 6.075 11.205 ;
        RECT 6.625 11.035 6.795 11.205 ;
        RECT 7.085 11.035 7.255 11.205 ;
        RECT 7.545 11.035 7.715 11.205 ;
        RECT 8.225 11.035 8.395 11.205 ;
        RECT 8.685 11.035 8.855 11.205 ;
        RECT 9.145 11.035 9.315 11.205 ;
        RECT 9.865 11.035 10.035 11.205 ;
        RECT 10.325 11.035 10.495 11.205 ;
        RECT 10.785 11.035 10.955 11.205 ;
        RECT 11.465 11.035 11.635 11.205 ;
        RECT 11.925 11.035 12.095 11.205 ;
        RECT 12.385 11.035 12.555 11.205 ;
        RECT 13.105 11.035 13.275 11.205 ;
        RECT 13.565 11.035 13.735 11.205 ;
        RECT 14.025 11.035 14.195 11.205 ;
        RECT 14.705 11.035 14.875 11.205 ;
        RECT 15.165 11.035 15.335 11.205 ;
        RECT 15.625 11.035 15.795 11.205 ;
        RECT 16.345 11.035 16.515 11.205 ;
        RECT 16.805 11.035 16.975 11.205 ;
        RECT 17.265 11.035 17.435 11.205 ;
        RECT 17.945 11.035 18.115 11.205 ;
        RECT 18.405 11.035 18.575 11.205 ;
        RECT 18.865 11.035 19.035 11.205 ;
        RECT 19.585 11.035 19.755 11.205 ;
        RECT 20.045 11.035 20.215 11.205 ;
        RECT 20.505 11.035 20.675 11.205 ;
        RECT 21.185 11.035 21.355 11.205 ;
        RECT 21.645 11.035 21.815 11.205 ;
        RECT 22.105 11.035 22.275 11.205 ;
        RECT 0.965 8.715 1.135 8.885 ;
        RECT 1.395 8.715 1.565 8.885 ;
        RECT 2.665 8.715 2.835 8.885 ;
        RECT 4.205 8.715 4.375 8.885 ;
        RECT 4.635 8.715 4.805 8.885 ;
        RECT 5.905 8.715 6.075 8.885 ;
        RECT 7.445 8.715 7.615 8.885 ;
        RECT 7.875 8.715 8.045 8.885 ;
        RECT 9.145 8.715 9.315 8.885 ;
        RECT 10.685 8.715 10.855 8.885 ;
        RECT 11.115 8.715 11.285 8.885 ;
        RECT 12.385 8.715 12.555 8.885 ;
        RECT 13.925 8.715 14.095 8.885 ;
        RECT 14.355 8.715 14.525 8.885 ;
        RECT 15.625 8.715 15.795 8.885 ;
        RECT 17.165 8.715 17.335 8.885 ;
        RECT 17.595 8.715 17.765 8.885 ;
        RECT 18.865 8.715 19.035 8.885 ;
        RECT 20.405 8.715 20.575 8.885 ;
        RECT 20.835 8.715 21.005 8.885 ;
        RECT 22.105 8.715 22.275 8.885 ;
        RECT 0.400 6.985 0.570 7.155 ;
        RECT 0.400 6.625 0.570 6.795 ;
        RECT 0.400 6.265 0.570 6.435 ;
        RECT 1.880 6.985 2.050 7.155 ;
        RECT 1.880 6.625 2.050 6.795 ;
        RECT 1.880 6.265 2.050 6.435 ;
        RECT 3.640 6.985 3.810 7.155 ;
        RECT 3.640 6.625 3.810 6.795 ;
        RECT 3.640 6.265 3.810 6.435 ;
        RECT 5.120 6.985 5.290 7.155 ;
        RECT 5.120 6.625 5.290 6.795 ;
        RECT 5.120 6.265 5.290 6.435 ;
        RECT 6.880 6.985 7.050 7.155 ;
        RECT 6.880 6.625 7.050 6.795 ;
        RECT 6.880 6.265 7.050 6.435 ;
        RECT 8.360 6.985 8.530 7.155 ;
        RECT 8.360 6.625 8.530 6.795 ;
        RECT 8.360 6.265 8.530 6.435 ;
        RECT 10.120 6.985 10.290 7.155 ;
        RECT 10.120 6.625 10.290 6.795 ;
        RECT 10.120 6.265 10.290 6.435 ;
        RECT 11.600 6.985 11.770 7.155 ;
        RECT 11.600 6.625 11.770 6.795 ;
        RECT 11.600 6.265 11.770 6.435 ;
        RECT 13.360 6.985 13.530 7.155 ;
        RECT 13.360 6.625 13.530 6.795 ;
        RECT 13.360 6.265 13.530 6.435 ;
        RECT 14.840 6.985 15.010 7.155 ;
        RECT 14.840 6.625 15.010 6.795 ;
        RECT 14.840 6.265 15.010 6.435 ;
        RECT 16.600 6.985 16.770 7.155 ;
        RECT 16.600 6.625 16.770 6.795 ;
        RECT 16.600 6.265 16.770 6.435 ;
        RECT 18.080 6.985 18.250 7.155 ;
        RECT 18.080 6.625 18.250 6.795 ;
        RECT 18.080 6.265 18.250 6.435 ;
        RECT 19.840 6.985 20.010 7.155 ;
        RECT 19.840 6.625 20.010 6.795 ;
        RECT 19.840 6.265 20.010 6.435 ;
        RECT 21.320 6.985 21.490 7.155 ;
        RECT 21.320 6.625 21.490 6.795 ;
        RECT 21.320 6.265 21.490 6.435 ;
        RECT 1.190 4.865 1.360 5.035 ;
        RECT 1.190 4.505 1.360 4.675 ;
        RECT 1.190 4.145 1.360 4.315 ;
        RECT 2.670 4.865 2.840 5.035 ;
        RECT 2.670 4.505 2.840 4.675 ;
        RECT 2.670 4.145 2.840 4.315 ;
        RECT 4.430 4.865 4.600 5.035 ;
        RECT 4.430 4.505 4.600 4.675 ;
        RECT 4.430 4.145 4.600 4.315 ;
        RECT 5.910 4.865 6.080 5.035 ;
        RECT 5.910 4.505 6.080 4.675 ;
        RECT 5.910 4.145 6.080 4.315 ;
        RECT 7.670 4.865 7.840 5.035 ;
        RECT 7.670 4.505 7.840 4.675 ;
        RECT 7.670 4.145 7.840 4.315 ;
        RECT 9.150 4.865 9.320 5.035 ;
        RECT 9.150 4.505 9.320 4.675 ;
        RECT 9.150 4.145 9.320 4.315 ;
        RECT 10.910 4.865 11.080 5.035 ;
        RECT 10.910 4.505 11.080 4.675 ;
        RECT 10.910 4.145 11.080 4.315 ;
        RECT 12.390 4.865 12.560 5.035 ;
        RECT 12.390 4.505 12.560 4.675 ;
        RECT 12.390 4.145 12.560 4.315 ;
        RECT 14.150 4.865 14.320 5.035 ;
        RECT 14.150 4.505 14.320 4.675 ;
        RECT 14.150 4.145 14.320 4.315 ;
        RECT 15.630 4.865 15.800 5.035 ;
        RECT 15.630 4.505 15.800 4.675 ;
        RECT 15.630 4.145 15.800 4.315 ;
        RECT 17.390 4.865 17.560 5.035 ;
        RECT 17.390 4.505 17.560 4.675 ;
        RECT 17.390 4.145 17.560 4.315 ;
        RECT 18.870 4.865 19.040 5.035 ;
        RECT 18.870 4.505 19.040 4.675 ;
        RECT 18.870 4.145 19.040 4.315 ;
        RECT 20.630 4.865 20.800 5.035 ;
        RECT 20.630 4.505 20.800 4.675 ;
        RECT 20.630 4.145 20.800 4.315 ;
        RECT 22.110 4.865 22.280 5.035 ;
        RECT 22.110 4.505 22.280 4.675 ;
        RECT 22.110 4.145 22.280 4.315 ;
        RECT 0.405 2.475 0.575 2.645 ;
        RECT 1.675 2.475 1.845 2.645 ;
        RECT 2.105 2.475 2.275 2.645 ;
        RECT 3.645 2.475 3.815 2.645 ;
        RECT 4.915 2.475 5.085 2.645 ;
        RECT 5.345 2.475 5.515 2.645 ;
        RECT 6.885 2.475 7.055 2.645 ;
        RECT 8.155 2.475 8.325 2.645 ;
        RECT 8.585 2.475 8.755 2.645 ;
        RECT 10.125 2.475 10.295 2.645 ;
        RECT 11.395 2.475 11.565 2.645 ;
        RECT 11.825 2.475 11.995 2.645 ;
        RECT 13.365 2.475 13.535 2.645 ;
        RECT 14.635 2.475 14.805 2.645 ;
        RECT 15.065 2.475 15.235 2.645 ;
        RECT 16.605 2.475 16.775 2.645 ;
        RECT 17.875 2.475 18.045 2.645 ;
        RECT 18.305 2.475 18.475 2.645 ;
        RECT 19.845 2.475 20.015 2.645 ;
        RECT 21.115 2.475 21.285 2.645 ;
        RECT 21.545 2.475 21.715 2.645 ;
        RECT 0.405 0.155 0.575 0.325 ;
        RECT 0.865 0.155 1.035 0.325 ;
        RECT 1.325 0.155 1.495 0.325 ;
        RECT 2.005 0.155 2.175 0.325 ;
        RECT 2.465 0.155 2.635 0.325 ;
        RECT 2.925 0.155 3.095 0.325 ;
        RECT 3.645 0.155 3.815 0.325 ;
        RECT 4.105 0.155 4.275 0.325 ;
        RECT 4.565 0.155 4.735 0.325 ;
        RECT 5.245 0.155 5.415 0.325 ;
        RECT 5.705 0.155 5.875 0.325 ;
        RECT 6.165 0.155 6.335 0.325 ;
        RECT 6.885 0.155 7.055 0.325 ;
        RECT 7.345 0.155 7.515 0.325 ;
        RECT 7.805 0.155 7.975 0.325 ;
        RECT 8.485 0.155 8.655 0.325 ;
        RECT 8.945 0.155 9.115 0.325 ;
        RECT 9.405 0.155 9.575 0.325 ;
        RECT 10.125 0.155 10.295 0.325 ;
        RECT 10.585 0.155 10.755 0.325 ;
        RECT 11.045 0.155 11.215 0.325 ;
        RECT 11.725 0.155 11.895 0.325 ;
        RECT 12.185 0.155 12.355 0.325 ;
        RECT 12.645 0.155 12.815 0.325 ;
        RECT 13.365 0.155 13.535 0.325 ;
        RECT 13.825 0.155 13.995 0.325 ;
        RECT 14.285 0.155 14.455 0.325 ;
        RECT 14.965 0.155 15.135 0.325 ;
        RECT 15.425 0.155 15.595 0.325 ;
        RECT 15.885 0.155 16.055 0.325 ;
        RECT 16.605 0.155 16.775 0.325 ;
        RECT 17.065 0.155 17.235 0.325 ;
        RECT 17.525 0.155 17.695 0.325 ;
        RECT 18.205 0.155 18.375 0.325 ;
        RECT 18.665 0.155 18.835 0.325 ;
        RECT 19.125 0.155 19.295 0.325 ;
        RECT 19.845 0.155 20.015 0.325 ;
        RECT 20.305 0.155 20.475 0.325 ;
        RECT 20.765 0.155 20.935 0.325 ;
        RECT 21.445 0.155 21.615 0.325 ;
        RECT 21.905 0.155 22.075 0.325 ;
        RECT 22.365 0.155 22.535 0.325 ;
      LAYER met1 ;
        RECT 0.000 10.880 22.680 11.360 ;
        RECT 0.000 8.670 22.680 9.040 ;
        RECT 0.370 7.010 0.600 7.400 ;
        RECT 1.850 7.010 2.080 7.400 ;
        RECT 3.610 7.010 3.840 7.400 ;
        RECT 5.090 7.010 5.320 7.400 ;
        RECT 6.850 7.010 7.080 7.400 ;
        RECT 8.330 7.010 8.560 7.400 ;
        RECT 10.090 7.010 10.320 7.400 ;
        RECT 11.570 7.010 11.800 7.400 ;
        RECT 13.330 7.010 13.560 7.400 ;
        RECT 14.810 7.010 15.040 7.400 ;
        RECT 16.570 7.010 16.800 7.400 ;
        RECT 18.050 7.010 18.280 7.400 ;
        RECT 19.810 7.010 20.040 7.400 ;
        RECT 21.290 7.010 21.520 7.400 ;
        RECT 0.280 6.750 0.600 7.010 ;
        RECT 1.760 6.750 2.080 7.010 ;
        RECT 3.520 6.750 3.840 7.010 ;
        RECT 5.000 6.750 5.320 7.010 ;
        RECT 6.760 6.750 7.080 7.010 ;
        RECT 8.240 6.750 8.560 7.010 ;
        RECT 10.000 6.750 10.320 7.010 ;
        RECT 11.480 6.750 11.800 7.010 ;
        RECT 13.240 6.750 13.560 7.010 ;
        RECT 14.720 6.750 15.040 7.010 ;
        RECT 16.480 6.750 16.800 7.010 ;
        RECT 17.960 6.750 18.280 7.010 ;
        RECT 19.720 6.750 20.040 7.010 ;
        RECT 21.200 6.750 21.520 7.010 ;
        RECT 0.370 6.140 0.600 6.750 ;
        RECT 1.850 6.140 2.080 6.750 ;
        RECT 3.610 6.140 3.840 6.750 ;
        RECT 5.090 6.140 5.320 6.750 ;
        RECT 6.850 6.140 7.080 6.750 ;
        RECT 8.330 6.140 8.560 6.750 ;
        RECT 10.090 6.140 10.320 6.750 ;
        RECT 11.570 6.140 11.800 6.750 ;
        RECT 13.330 6.140 13.560 6.750 ;
        RECT 14.810 6.140 15.040 6.750 ;
        RECT 16.570 6.140 16.800 6.750 ;
        RECT 18.050 6.140 18.280 6.750 ;
        RECT 19.810 6.140 20.040 6.750 ;
        RECT 21.290 6.140 21.520 6.750 ;
        RECT 1.160 4.510 1.390 5.160 ;
        RECT 2.640 4.510 2.870 5.160 ;
        RECT 4.400 4.510 4.630 5.160 ;
        RECT 5.880 4.510 6.110 5.160 ;
        RECT 7.640 4.510 7.870 5.160 ;
        RECT 9.120 4.510 9.350 5.160 ;
        RECT 10.880 4.510 11.110 5.160 ;
        RECT 12.360 4.510 12.590 5.160 ;
        RECT 14.120 4.510 14.350 5.160 ;
        RECT 15.600 4.510 15.830 5.160 ;
        RECT 17.360 4.510 17.590 5.160 ;
        RECT 18.840 4.510 19.070 5.160 ;
        RECT 20.600 4.510 20.830 5.160 ;
        RECT 22.080 4.510 22.310 5.160 ;
        RECT 1.160 4.250 1.480 4.510 ;
        RECT 2.640 4.250 2.960 4.510 ;
        RECT 4.400 4.250 4.720 4.510 ;
        RECT 5.880 4.250 6.200 4.510 ;
        RECT 7.640 4.250 7.960 4.510 ;
        RECT 9.120 4.250 9.440 4.510 ;
        RECT 10.880 4.250 11.200 4.510 ;
        RECT 12.360 4.250 12.680 4.510 ;
        RECT 14.120 4.250 14.440 4.510 ;
        RECT 15.600 4.250 15.920 4.510 ;
        RECT 17.360 4.250 17.680 4.510 ;
        RECT 18.840 4.250 19.160 4.510 ;
        RECT 20.600 4.250 20.920 4.510 ;
        RECT 22.080 4.250 22.400 4.510 ;
        RECT 1.160 3.900 1.390 4.250 ;
        RECT 2.640 3.900 2.870 4.250 ;
        RECT 4.400 3.900 4.630 4.250 ;
        RECT 5.880 3.900 6.110 4.250 ;
        RECT 7.640 3.900 7.870 4.250 ;
        RECT 9.120 3.900 9.350 4.250 ;
        RECT 10.880 3.900 11.110 4.250 ;
        RECT 12.360 3.900 12.590 4.250 ;
        RECT 14.120 3.900 14.350 4.250 ;
        RECT 15.600 3.900 15.830 4.250 ;
        RECT 17.360 3.900 17.590 4.250 ;
        RECT 18.840 3.900 19.070 4.250 ;
        RECT 20.600 3.900 20.830 4.250 ;
        RECT 22.080 3.900 22.310 4.250 ;
        RECT 0.000 2.320 22.680 2.690 ;
        RECT 0.000 0.000 22.680 0.480 ;
  END
END rram_28
END LIBRARY

