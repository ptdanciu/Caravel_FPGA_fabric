VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS
MACRO test_lut_inst
  FOREIGN test_lut_inst 0 0 ;
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 352.05 BY 202 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      VIA 334.8 195.88 via4_1600x1600 ;
      VIA 314.6 195.88 via4_1600x1600 ;
      VIA 294.4 195.88 via4_1600x1600 ;
      VIA 274.2 195.88 via4_1600x1600 ;
      VIA 254 195.88 via4_1600x1600 ;
      VIA 233.8 195.88 via4_1600x1600 ;
      VIA 213.6 195.88 via4_1600x1600 ;
      VIA 193.4 195.88 via4_1600x1600 ;
      VIA 173.2 195.88 via4_1600x1600 ;
      VIA 153 195.88 via4_1600x1600 ;
      VIA 132.8 195.88 via4_1600x1600 ;
      VIA 112.6 195.88 via4_1600x1600 ;
      VIA 92.4 195.88 via4_1600x1600 ;
      VIA 72.2 195.88 via4_1600x1600 ;
      VIA 52 195.88 via4_1600x1600 ;
      VIA 31.8 195.88 via4_1600x1600 ;
      VIA 11.6 195.88 via4_1600x1600 ;
      VIA 334.8 175.68 via4_1600x1600 ;
      VIA 314.6 175.68 via4_1600x1600 ;
      VIA 294.4 175.68 via4_1600x1600 ;
      VIA 274.2 175.68 via4_1600x1600 ;
      VIA 254 175.68 via4_1600x1600 ;
      VIA 233.8 175.68 via4_1600x1600 ;
      VIA 213.6 175.68 via4_1600x1600 ;
      VIA 193.4 175.68 via4_1600x1600 ;
      VIA 173.2 175.68 via4_1600x1600 ;
      VIA 153 175.68 via4_1600x1600 ;
      VIA 132.8 175.68 via4_1600x1600 ;
      VIA 112.6 175.68 via4_1600x1600 ;
      VIA 92.4 175.68 via4_1600x1600 ;
      VIA 72.2 175.68 via4_1600x1600 ;
      VIA 52 175.68 via4_1600x1600 ;
      VIA 31.8 175.68 via4_1600x1600 ;
      VIA 11.6 175.68 via4_1600x1600 ;
      VIA 334.8 155.48 via4_1600x1600 ;
      VIA 314.6 155.48 via4_1600x1600 ;
      VIA 294.4 155.48 via4_1600x1600 ;
      VIA 274.2 155.48 via4_1600x1600 ;
      VIA 254 155.48 via4_1600x1600 ;
      VIA 233.8 155.48 via4_1600x1600 ;
      VIA 213.6 155.48 via4_1600x1600 ;
      VIA 193.4 155.48 via4_1600x1600 ;
      VIA 173.2 155.48 via4_1600x1600 ;
      VIA 153 155.48 via4_1600x1600 ;
      VIA 132.8 155.48 via4_1600x1600 ;
      VIA 112.6 155.48 via4_1600x1600 ;
      VIA 92.4 155.48 via4_1600x1600 ;
      VIA 72.2 155.48 via4_1600x1600 ;
      VIA 52 155.48 via4_1600x1600 ;
      VIA 31.8 155.48 via4_1600x1600 ;
      VIA 11.6 155.48 via4_1600x1600 ;
      VIA 334.8 135.28 via4_1600x1600 ;
      VIA 314.6 135.28 via4_1600x1600 ;
      VIA 294.4 135.28 via4_1600x1600 ;
      VIA 274.2 135.28 via4_1600x1600 ;
      VIA 254 135.28 via4_1600x1600 ;
      VIA 233.8 135.28 via4_1600x1600 ;
      VIA 213.6 135.28 via4_1600x1600 ;
      VIA 193.4 135.28 via4_1600x1600 ;
      VIA 173.2 135.28 via4_1600x1600 ;
      VIA 153 135.28 via4_1600x1600 ;
      VIA 132.8 135.28 via4_1600x1600 ;
      VIA 112.6 135.28 via4_1600x1600 ;
      VIA 92.4 135.28 via4_1600x1600 ;
      VIA 72.2 135.28 via4_1600x1600 ;
      VIA 52 135.28 via4_1600x1600 ;
      VIA 31.8 135.28 via4_1600x1600 ;
      VIA 11.6 135.28 via4_1600x1600 ;
      VIA 334.8 115.08 via4_1600x1600 ;
      VIA 314.6 115.08 via4_1600x1600 ;
      VIA 294.4 115.08 via4_1600x1600 ;
      VIA 274.2 115.08 via4_1600x1600 ;
      VIA 254 115.08 via4_1600x1600 ;
      VIA 233.8 115.08 via4_1600x1600 ;
      VIA 213.6 115.08 via4_1600x1600 ;
      VIA 193.4 115.08 via4_1600x1600 ;
      VIA 173.2 115.08 via4_1600x1600 ;
      VIA 153 115.08 via4_1600x1600 ;
      VIA 132.8 115.08 via4_1600x1600 ;
      VIA 112.6 115.08 via4_1600x1600 ;
      VIA 92.4 115.08 via4_1600x1600 ;
      VIA 72.2 115.08 via4_1600x1600 ;
      VIA 52 115.08 via4_1600x1600 ;
      VIA 31.8 115.08 via4_1600x1600 ;
      VIA 11.6 115.08 via4_1600x1600 ;
      VIA 334.8 94.88 via4_1600x1600 ;
      VIA 314.6 94.88 via4_1600x1600 ;
      VIA 294.4 94.88 via4_1600x1600 ;
      VIA 274.2 94.88 via4_1600x1600 ;
      VIA 254 94.88 via4_1600x1600 ;
      VIA 233.8 94.88 via4_1600x1600 ;
      VIA 213.6 94.88 via4_1600x1600 ;
      VIA 193.4 94.88 via4_1600x1600 ;
      VIA 173.2 94.88 via4_1600x1600 ;
      VIA 153 94.88 via4_1600x1600 ;
      VIA 132.8 94.88 via4_1600x1600 ;
      VIA 112.6 94.88 via4_1600x1600 ;
      VIA 92.4 94.88 via4_1600x1600 ;
      VIA 72.2 94.88 via4_1600x1600 ;
      VIA 52 94.88 via4_1600x1600 ;
      VIA 31.8 94.88 via4_1600x1600 ;
      VIA 11.6 94.88 via4_1600x1600 ;
      VIA 334.8 74.68 via4_1600x1600 ;
      VIA 314.6 74.68 via4_1600x1600 ;
      VIA 294.4 74.68 via4_1600x1600 ;
      VIA 274.2 74.68 via4_1600x1600 ;
      VIA 254 74.68 via4_1600x1600 ;
      VIA 233.8 74.68 via4_1600x1600 ;
      VIA 213.6 74.68 via4_1600x1600 ;
      VIA 193.4 74.68 via4_1600x1600 ;
      VIA 173.2 74.68 via4_1600x1600 ;
      VIA 153 74.68 via4_1600x1600 ;
      VIA 132.8 74.68 via4_1600x1600 ;
      VIA 112.6 74.68 via4_1600x1600 ;
      VIA 92.4 74.68 via4_1600x1600 ;
      VIA 72.2 74.68 via4_1600x1600 ;
      VIA 52 74.68 via4_1600x1600 ;
      VIA 31.8 74.68 via4_1600x1600 ;
      VIA 11.6 74.68 via4_1600x1600 ;
      VIA 334.8 54.48 via4_1600x1600 ;
      VIA 314.6 54.48 via4_1600x1600 ;
      VIA 294.4 54.48 via4_1600x1600 ;
      VIA 274.2 54.48 via4_1600x1600 ;
      VIA 254 54.48 via4_1600x1600 ;
      VIA 233.8 54.48 via4_1600x1600 ;
      VIA 213.6 54.48 via4_1600x1600 ;
      VIA 193.4 54.48 via4_1600x1600 ;
      VIA 173.2 54.48 via4_1600x1600 ;
      VIA 153 54.48 via4_1600x1600 ;
      VIA 132.8 54.48 via4_1600x1600 ;
      VIA 112.6 54.48 via4_1600x1600 ;
      VIA 92.4 54.48 via4_1600x1600 ;
      VIA 72.2 54.48 via4_1600x1600 ;
      VIA 52 54.48 via4_1600x1600 ;
      VIA 31.8 54.48 via4_1600x1600 ;
      VIA 11.6 54.48 via4_1600x1600 ;
      VIA 334.8 34.28 via4_1600x1600 ;
      VIA 314.6 34.28 via4_1600x1600 ;
      VIA 294.4 34.28 via4_1600x1600 ;
      VIA 274.2 34.28 via4_1600x1600 ;
      VIA 254 34.28 via4_1600x1600 ;
      VIA 233.8 34.28 via4_1600x1600 ;
      VIA 213.6 34.28 via4_1600x1600 ;
      VIA 193.4 34.28 via4_1600x1600 ;
      VIA 173.2 34.28 via4_1600x1600 ;
      VIA 153 34.28 via4_1600x1600 ;
      VIA 132.8 34.28 via4_1600x1600 ;
      VIA 112.6 34.28 via4_1600x1600 ;
      VIA 92.4 34.28 via4_1600x1600 ;
      VIA 72.2 34.28 via4_1600x1600 ;
      VIA 52 34.28 via4_1600x1600 ;
      VIA 31.8 34.28 via4_1600x1600 ;
      VIA 11.6 34.28 via4_1600x1600 ;
      VIA 334.8 14.08 via4_1600x1600 ;
      VIA 314.6 14.08 via4_1600x1600 ;
      VIA 294.4 14.08 via4_1600x1600 ;
      VIA 274.2 14.08 via4_1600x1600 ;
      VIA 254 14.08 via4_1600x1600 ;
      VIA 233.8 14.08 via4_1600x1600 ;
      VIA 213.6 14.08 via4_1600x1600 ;
      VIA 193.4 14.08 via4_1600x1600 ;
      VIA 173.2 14.08 via4_1600x1600 ;
      VIA 153 14.08 via4_1600x1600 ;
      VIA 132.8 14.08 via4_1600x1600 ;
      VIA 112.6 14.08 via4_1600x1600 ;
      VIA 92.4 14.08 via4_1600x1600 ;
      VIA 72.2 14.08 via4_1600x1600 ;
      VIA 52 14.08 via4_1600x1600 ;
      VIA 31.8 14.08 via4_1600x1600 ;
      VIA 11.6 14.08 via4_1600x1600 ;
      VIA 334.8 195.84 via3_1600x480 ;
      VIA 334.8 195.84 via2_1600x480 ;
      VIA 334.8 195.84 via_1600x480 ;
      VIA 314.6 195.84 via3_1600x480 ;
      VIA 314.6 195.84 via2_1600x480 ;
      VIA 314.6 195.84 via_1600x480 ;
      VIA 294.4 195.84 via3_1600x480 ;
      VIA 294.4 195.84 via2_1600x480 ;
      VIA 294.4 195.84 via_1600x480 ;
      VIA 274.2 195.84 via3_1600x480 ;
      VIA 274.2 195.84 via2_1600x480 ;
      VIA 274.2 195.84 via_1600x480 ;
      VIA 254 195.84 via3_1600x480 ;
      VIA 254 195.84 via2_1600x480 ;
      VIA 254 195.84 via_1600x480 ;
      VIA 233.8 195.84 via3_1600x480 ;
      VIA 233.8 195.84 via2_1600x480 ;
      VIA 233.8 195.84 via_1600x480 ;
      VIA 213.6 195.84 via3_1600x480 ;
      VIA 213.6 195.84 via2_1600x480 ;
      VIA 213.6 195.84 via_1600x480 ;
      VIA 193.4 195.84 via3_1600x480 ;
      VIA 193.4 195.84 via2_1600x480 ;
      VIA 193.4 195.84 via_1600x480 ;
      VIA 173.2 195.84 via3_1600x480 ;
      VIA 173.2 195.84 via2_1600x480 ;
      VIA 173.2 195.84 via_1600x480 ;
      VIA 153 195.84 via3_1600x480 ;
      VIA 153 195.84 via2_1600x480 ;
      VIA 153 195.84 via_1600x480 ;
      VIA 132.8 195.84 via3_1600x480 ;
      VIA 132.8 195.84 via2_1600x480 ;
      VIA 132.8 195.84 via_1600x480 ;
      VIA 112.6 195.84 via3_1600x480 ;
      VIA 112.6 195.84 via2_1600x480 ;
      VIA 112.6 195.84 via_1600x480 ;
      VIA 92.4 195.84 via3_1600x480 ;
      VIA 92.4 195.84 via2_1600x480 ;
      VIA 92.4 195.84 via_1600x480 ;
      VIA 72.2 195.84 via3_1600x480 ;
      VIA 72.2 195.84 via2_1600x480 ;
      VIA 72.2 195.84 via_1600x480 ;
      VIA 52 195.84 via3_1600x480 ;
      VIA 52 195.84 via2_1600x480 ;
      VIA 52 195.84 via_1600x480 ;
      VIA 31.8 195.84 via3_1600x480 ;
      VIA 31.8 195.84 via2_1600x480 ;
      VIA 31.8 195.84 via_1600x480 ;
      VIA 11.6 195.84 via3_1600x480 ;
      VIA 11.6 195.84 via2_1600x480 ;
      VIA 11.6 195.84 via_1600x480 ;
      VIA 334.8 190.4 via3_1600x480 ;
      VIA 334.8 190.4 via2_1600x480 ;
      VIA 334.8 190.4 via_1600x480 ;
      VIA 314.6 190.4 via3_1600x480 ;
      VIA 314.6 190.4 via2_1600x480 ;
      VIA 314.6 190.4 via_1600x480 ;
      VIA 294.4 190.4 via3_1600x480 ;
      VIA 294.4 190.4 via2_1600x480 ;
      VIA 294.4 190.4 via_1600x480 ;
      VIA 274.2 190.4 via3_1600x480 ;
      VIA 274.2 190.4 via2_1600x480 ;
      VIA 274.2 190.4 via_1600x480 ;
      VIA 254 190.4 via3_1600x480 ;
      VIA 254 190.4 via2_1600x480 ;
      VIA 254 190.4 via_1600x480 ;
      VIA 233.8 190.4 via3_1600x480 ;
      VIA 233.8 190.4 via2_1600x480 ;
      VIA 233.8 190.4 via_1600x480 ;
      VIA 213.6 190.4 via3_1600x480 ;
      VIA 213.6 190.4 via2_1600x480 ;
      VIA 213.6 190.4 via_1600x480 ;
      VIA 193.4 190.4 via3_1600x480 ;
      VIA 193.4 190.4 via2_1600x480 ;
      VIA 193.4 190.4 via_1600x480 ;
      VIA 173.2 190.4 via3_1600x480 ;
      VIA 173.2 190.4 via2_1600x480 ;
      VIA 173.2 190.4 via_1600x480 ;
      VIA 153 190.4 via3_1600x480 ;
      VIA 153 190.4 via2_1600x480 ;
      VIA 153 190.4 via_1600x480 ;
      VIA 132.8 190.4 via3_1600x480 ;
      VIA 132.8 190.4 via2_1600x480 ;
      VIA 132.8 190.4 via_1600x480 ;
      VIA 112.6 190.4 via3_1600x480 ;
      VIA 112.6 190.4 via2_1600x480 ;
      VIA 112.6 190.4 via_1600x480 ;
      VIA 92.4 190.4 via3_1600x480 ;
      VIA 92.4 190.4 via2_1600x480 ;
      VIA 92.4 190.4 via_1600x480 ;
      VIA 72.2 190.4 via3_1600x480 ;
      VIA 72.2 190.4 via2_1600x480 ;
      VIA 72.2 190.4 via_1600x480 ;
      VIA 52 190.4 via3_1600x480 ;
      VIA 52 190.4 via2_1600x480 ;
      VIA 52 190.4 via_1600x480 ;
      VIA 31.8 190.4 via3_1600x480 ;
      VIA 31.8 190.4 via2_1600x480 ;
      VIA 31.8 190.4 via_1600x480 ;
      VIA 11.6 190.4 via3_1600x480 ;
      VIA 11.6 190.4 via2_1600x480 ;
      VIA 11.6 190.4 via_1600x480 ;
      VIA 334.8 184.96 via3_1600x480 ;
      VIA 334.8 184.96 via2_1600x480 ;
      VIA 334.8 184.96 via_1600x480 ;
      VIA 314.6 184.96 via3_1600x480 ;
      VIA 314.6 184.96 via2_1600x480 ;
      VIA 314.6 184.96 via_1600x480 ;
      VIA 294.4 184.96 via3_1600x480 ;
      VIA 294.4 184.96 via2_1600x480 ;
      VIA 294.4 184.96 via_1600x480 ;
      VIA 274.2 184.96 via3_1600x480 ;
      VIA 274.2 184.96 via2_1600x480 ;
      VIA 274.2 184.96 via_1600x480 ;
      VIA 254 184.96 via3_1600x480 ;
      VIA 254 184.96 via2_1600x480 ;
      VIA 254 184.96 via_1600x480 ;
      VIA 233.8 184.96 via3_1600x480 ;
      VIA 233.8 184.96 via2_1600x480 ;
      VIA 233.8 184.96 via_1600x480 ;
      VIA 213.6 184.96 via3_1600x480 ;
      VIA 213.6 184.96 via2_1600x480 ;
      VIA 213.6 184.96 via_1600x480 ;
      VIA 193.4 184.96 via3_1600x480 ;
      VIA 193.4 184.96 via2_1600x480 ;
      VIA 193.4 184.96 via_1600x480 ;
      VIA 173.2 184.96 via3_1600x480 ;
      VIA 173.2 184.96 via2_1600x480 ;
      VIA 173.2 184.96 via_1600x480 ;
      VIA 153 184.96 via3_1600x480 ;
      VIA 153 184.96 via2_1600x480 ;
      VIA 153 184.96 via_1600x480 ;
      VIA 132.8 184.96 via3_1600x480 ;
      VIA 132.8 184.96 via2_1600x480 ;
      VIA 132.8 184.96 via_1600x480 ;
      VIA 112.6 184.96 via3_1600x480 ;
      VIA 112.6 184.96 via2_1600x480 ;
      VIA 112.6 184.96 via_1600x480 ;
      VIA 92.4 184.96 via3_1600x480 ;
      VIA 92.4 184.96 via2_1600x480 ;
      VIA 92.4 184.96 via_1600x480 ;
      VIA 72.2 184.96 via3_1600x480 ;
      VIA 72.2 184.96 via2_1600x480 ;
      VIA 72.2 184.96 via_1600x480 ;
      VIA 52 184.96 via3_1600x480 ;
      VIA 52 184.96 via2_1600x480 ;
      VIA 52 184.96 via_1600x480 ;
      VIA 31.8 184.96 via3_1600x480 ;
      VIA 31.8 184.96 via2_1600x480 ;
      VIA 31.8 184.96 via_1600x480 ;
      VIA 11.6 184.96 via3_1600x480 ;
      VIA 11.6 184.96 via2_1600x480 ;
      VIA 11.6 184.96 via_1600x480 ;
      VIA 334.8 179.52 via3_1600x480 ;
      VIA 334.8 179.52 via2_1600x480 ;
      VIA 334.8 179.52 via_1600x480 ;
      VIA 314.6 179.52 via3_1600x480 ;
      VIA 314.6 179.52 via2_1600x480 ;
      VIA 314.6 179.52 via_1600x480 ;
      VIA 294.4 179.52 via3_1600x480 ;
      VIA 294.4 179.52 via2_1600x480 ;
      VIA 294.4 179.52 via_1600x480 ;
      VIA 274.2 179.52 via3_1600x480 ;
      VIA 274.2 179.52 via2_1600x480 ;
      VIA 274.2 179.52 via_1600x480 ;
      VIA 254 179.52 via3_1600x480 ;
      VIA 254 179.52 via2_1600x480 ;
      VIA 254 179.52 via_1600x480 ;
      VIA 233.8 179.52 via3_1600x480 ;
      VIA 233.8 179.52 via2_1600x480 ;
      VIA 233.8 179.52 via_1600x480 ;
      VIA 213.6 179.52 via3_1600x480 ;
      VIA 213.6 179.52 via2_1600x480 ;
      VIA 213.6 179.52 via_1600x480 ;
      VIA 193.4 179.52 via3_1600x480 ;
      VIA 193.4 179.52 via2_1600x480 ;
      VIA 193.4 179.52 via_1600x480 ;
      VIA 173.2 179.52 via3_1600x480 ;
      VIA 173.2 179.52 via2_1600x480 ;
      VIA 173.2 179.52 via_1600x480 ;
      VIA 153 179.52 via3_1600x480 ;
      VIA 153 179.52 via2_1600x480 ;
      VIA 153 179.52 via_1600x480 ;
      VIA 132.8 179.52 via3_1600x480 ;
      VIA 132.8 179.52 via2_1600x480 ;
      VIA 132.8 179.52 via_1600x480 ;
      VIA 112.6 179.52 via3_1600x480 ;
      VIA 112.6 179.52 via2_1600x480 ;
      VIA 112.6 179.52 via_1600x480 ;
      VIA 92.4 179.52 via3_1600x480 ;
      VIA 92.4 179.52 via2_1600x480 ;
      VIA 92.4 179.52 via_1600x480 ;
      VIA 72.2 179.52 via3_1600x480 ;
      VIA 72.2 179.52 via2_1600x480 ;
      VIA 72.2 179.52 via_1600x480 ;
      VIA 52 179.52 via3_1600x480 ;
      VIA 52 179.52 via2_1600x480 ;
      VIA 52 179.52 via_1600x480 ;
      VIA 31.8 179.52 via3_1600x480 ;
      VIA 31.8 179.52 via2_1600x480 ;
      VIA 31.8 179.52 via_1600x480 ;
      VIA 11.6 179.52 via3_1600x480 ;
      VIA 11.6 179.52 via2_1600x480 ;
      VIA 11.6 179.52 via_1600x480 ;
      VIA 334.8 174.08 via3_1600x480 ;
      VIA 334.8 174.08 via2_1600x480 ;
      VIA 334.8 174.08 via_1600x480 ;
      VIA 314.6 174.08 via3_1600x480 ;
      VIA 314.6 174.08 via2_1600x480 ;
      VIA 314.6 174.08 via_1600x480 ;
      VIA 294.4 174.08 via3_1600x480 ;
      VIA 294.4 174.08 via2_1600x480 ;
      VIA 294.4 174.08 via_1600x480 ;
      VIA 274.2 174.08 via3_1600x480 ;
      VIA 274.2 174.08 via2_1600x480 ;
      VIA 274.2 174.08 via_1600x480 ;
      VIA 254 174.08 via3_1600x480 ;
      VIA 254 174.08 via2_1600x480 ;
      VIA 254 174.08 via_1600x480 ;
      VIA 233.8 174.08 via3_1600x480 ;
      VIA 233.8 174.08 via2_1600x480 ;
      VIA 233.8 174.08 via_1600x480 ;
      VIA 213.6 174.08 via3_1600x480 ;
      VIA 213.6 174.08 via2_1600x480 ;
      VIA 213.6 174.08 via_1600x480 ;
      VIA 193.4 174.08 via3_1600x480 ;
      VIA 193.4 174.08 via2_1600x480 ;
      VIA 193.4 174.08 via_1600x480 ;
      VIA 173.2 174.08 via3_1600x480 ;
      VIA 173.2 174.08 via2_1600x480 ;
      VIA 173.2 174.08 via_1600x480 ;
      VIA 153 174.08 via3_1600x480 ;
      VIA 153 174.08 via2_1600x480 ;
      VIA 153 174.08 via_1600x480 ;
      VIA 132.8 174.08 via3_1600x480 ;
      VIA 132.8 174.08 via2_1600x480 ;
      VIA 132.8 174.08 via_1600x480 ;
      VIA 112.6 174.08 via3_1600x480 ;
      VIA 112.6 174.08 via2_1600x480 ;
      VIA 112.6 174.08 via_1600x480 ;
      VIA 92.4 174.08 via3_1600x480 ;
      VIA 92.4 174.08 via2_1600x480 ;
      VIA 92.4 174.08 via_1600x480 ;
      VIA 72.2 174.08 via3_1600x480 ;
      VIA 72.2 174.08 via2_1600x480 ;
      VIA 72.2 174.08 via_1600x480 ;
      VIA 52 174.08 via3_1600x480 ;
      VIA 52 174.08 via2_1600x480 ;
      VIA 52 174.08 via_1600x480 ;
      VIA 31.8 174.08 via3_1600x480 ;
      VIA 31.8 174.08 via2_1600x480 ;
      VIA 31.8 174.08 via_1600x480 ;
      VIA 11.6 174.08 via3_1600x480 ;
      VIA 11.6 174.08 via2_1600x480 ;
      VIA 11.6 174.08 via_1600x480 ;
      VIA 334.8 168.64 via3_1600x480 ;
      VIA 334.8 168.64 via2_1600x480 ;
      VIA 334.8 168.64 via_1600x480 ;
      VIA 314.6 168.64 via3_1600x480 ;
      VIA 314.6 168.64 via2_1600x480 ;
      VIA 314.6 168.64 via_1600x480 ;
      VIA 294.4 168.64 via3_1600x480 ;
      VIA 294.4 168.64 via2_1600x480 ;
      VIA 294.4 168.64 via_1600x480 ;
      VIA 274.2 168.64 via3_1600x480 ;
      VIA 274.2 168.64 via2_1600x480 ;
      VIA 274.2 168.64 via_1600x480 ;
      VIA 254 168.64 via3_1600x480 ;
      VIA 254 168.64 via2_1600x480 ;
      VIA 254 168.64 via_1600x480 ;
      VIA 233.8 168.64 via3_1600x480 ;
      VIA 233.8 168.64 via2_1600x480 ;
      VIA 233.8 168.64 via_1600x480 ;
      VIA 213.6 168.64 via3_1600x480 ;
      VIA 213.6 168.64 via2_1600x480 ;
      VIA 213.6 168.64 via_1600x480 ;
      VIA 193.4 168.64 via3_1600x480 ;
      VIA 193.4 168.64 via2_1600x480 ;
      VIA 193.4 168.64 via_1600x480 ;
      VIA 173.2 168.64 via3_1600x480 ;
      VIA 173.2 168.64 via2_1600x480 ;
      VIA 173.2 168.64 via_1600x480 ;
      VIA 153 168.64 via3_1600x480 ;
      VIA 153 168.64 via2_1600x480 ;
      VIA 153 168.64 via_1600x480 ;
      VIA 132.8 168.64 via3_1600x480 ;
      VIA 132.8 168.64 via2_1600x480 ;
      VIA 132.8 168.64 via_1600x480 ;
      VIA 112.6 168.64 via3_1600x480 ;
      VIA 112.6 168.64 via2_1600x480 ;
      VIA 112.6 168.64 via_1600x480 ;
      VIA 92.4 168.64 via3_1600x480 ;
      VIA 92.4 168.64 via2_1600x480 ;
      VIA 92.4 168.64 via_1600x480 ;
      VIA 72.2 168.64 via3_1600x480 ;
      VIA 72.2 168.64 via2_1600x480 ;
      VIA 72.2 168.64 via_1600x480 ;
      VIA 52 168.64 via3_1600x480 ;
      VIA 52 168.64 via2_1600x480 ;
      VIA 52 168.64 via_1600x480 ;
      VIA 31.8 168.64 via3_1600x480 ;
      VIA 31.8 168.64 via2_1600x480 ;
      VIA 31.8 168.64 via_1600x480 ;
      VIA 11.6 168.64 via3_1600x480 ;
      VIA 11.6 168.64 via2_1600x480 ;
      VIA 11.6 168.64 via_1600x480 ;
      VIA 334.8 163.2 via3_1600x480 ;
      VIA 334.8 163.2 via2_1600x480 ;
      VIA 334.8 163.2 via_1600x480 ;
      VIA 314.6 163.2 via3_1600x480 ;
      VIA 314.6 163.2 via2_1600x480 ;
      VIA 314.6 163.2 via_1600x480 ;
      VIA 294.4 163.2 via3_1600x480 ;
      VIA 294.4 163.2 via2_1600x480 ;
      VIA 294.4 163.2 via_1600x480 ;
      VIA 274.2 163.2 via3_1600x480 ;
      VIA 274.2 163.2 via2_1600x480 ;
      VIA 274.2 163.2 via_1600x480 ;
      VIA 254 163.2 via3_1600x480 ;
      VIA 254 163.2 via2_1600x480 ;
      VIA 254 163.2 via_1600x480 ;
      VIA 233.8 163.2 via3_1600x480 ;
      VIA 233.8 163.2 via2_1600x480 ;
      VIA 233.8 163.2 via_1600x480 ;
      VIA 213.6 163.2 via3_1600x480 ;
      VIA 213.6 163.2 via2_1600x480 ;
      VIA 213.6 163.2 via_1600x480 ;
      VIA 193.4 163.2 via3_1600x480 ;
      VIA 193.4 163.2 via2_1600x480 ;
      VIA 193.4 163.2 via_1600x480 ;
      VIA 173.2 163.2 via3_1600x480 ;
      VIA 173.2 163.2 via2_1600x480 ;
      VIA 173.2 163.2 via_1600x480 ;
      VIA 153 163.2 via3_1600x480 ;
      VIA 153 163.2 via2_1600x480 ;
      VIA 153 163.2 via_1600x480 ;
      VIA 132.8 163.2 via3_1600x480 ;
      VIA 132.8 163.2 via2_1600x480 ;
      VIA 132.8 163.2 via_1600x480 ;
      VIA 112.6 163.2 via3_1600x480 ;
      VIA 112.6 163.2 via2_1600x480 ;
      VIA 112.6 163.2 via_1600x480 ;
      VIA 92.4 163.2 via3_1600x480 ;
      VIA 92.4 163.2 via2_1600x480 ;
      VIA 92.4 163.2 via_1600x480 ;
      VIA 72.2 163.2 via3_1600x480 ;
      VIA 72.2 163.2 via2_1600x480 ;
      VIA 72.2 163.2 via_1600x480 ;
      VIA 52 163.2 via3_1600x480 ;
      VIA 52 163.2 via2_1600x480 ;
      VIA 52 163.2 via_1600x480 ;
      VIA 31.8 163.2 via3_1600x480 ;
      VIA 31.8 163.2 via2_1600x480 ;
      VIA 31.8 163.2 via_1600x480 ;
      VIA 11.6 163.2 via3_1600x480 ;
      VIA 11.6 163.2 via2_1600x480 ;
      VIA 11.6 163.2 via_1600x480 ;
      VIA 334.8 157.76 via3_1600x480 ;
      VIA 334.8 157.76 via2_1600x480 ;
      VIA 334.8 157.76 via_1600x480 ;
      VIA 314.6 157.76 via3_1600x480 ;
      VIA 314.6 157.76 via2_1600x480 ;
      VIA 314.6 157.76 via_1600x480 ;
      VIA 294.4 157.76 via3_1600x480 ;
      VIA 294.4 157.76 via2_1600x480 ;
      VIA 294.4 157.76 via_1600x480 ;
      VIA 274.2 157.76 via3_1600x480 ;
      VIA 274.2 157.76 via2_1600x480 ;
      VIA 274.2 157.76 via_1600x480 ;
      VIA 254 157.76 via3_1600x480 ;
      VIA 254 157.76 via2_1600x480 ;
      VIA 254 157.76 via_1600x480 ;
      VIA 233.8 157.76 via3_1600x480 ;
      VIA 233.8 157.76 via2_1600x480 ;
      VIA 233.8 157.76 via_1600x480 ;
      VIA 213.6 157.76 via3_1600x480 ;
      VIA 213.6 157.76 via2_1600x480 ;
      VIA 213.6 157.76 via_1600x480 ;
      VIA 193.4 157.76 via3_1600x480 ;
      VIA 193.4 157.76 via2_1600x480 ;
      VIA 193.4 157.76 via_1600x480 ;
      VIA 173.2 157.76 via3_1600x480 ;
      VIA 173.2 157.76 via2_1600x480 ;
      VIA 173.2 157.76 via_1600x480 ;
      VIA 153 157.76 via3_1600x480 ;
      VIA 153 157.76 via2_1600x480 ;
      VIA 153 157.76 via_1600x480 ;
      VIA 132.8 157.76 via3_1600x480 ;
      VIA 132.8 157.76 via2_1600x480 ;
      VIA 132.8 157.76 via_1600x480 ;
      VIA 112.6 157.76 via3_1600x480 ;
      VIA 112.6 157.76 via2_1600x480 ;
      VIA 112.6 157.76 via_1600x480 ;
      VIA 92.4 157.76 via3_1600x480 ;
      VIA 92.4 157.76 via2_1600x480 ;
      VIA 92.4 157.76 via_1600x480 ;
      VIA 72.2 157.76 via3_1600x480 ;
      VIA 72.2 157.76 via2_1600x480 ;
      VIA 72.2 157.76 via_1600x480 ;
      VIA 52 157.76 via3_1600x480 ;
      VIA 52 157.76 via2_1600x480 ;
      VIA 52 157.76 via_1600x480 ;
      VIA 31.8 157.76 via3_1600x480 ;
      VIA 31.8 157.76 via2_1600x480 ;
      VIA 31.8 157.76 via_1600x480 ;
      VIA 11.6 157.76 via3_1600x480 ;
      VIA 11.6 157.76 via2_1600x480 ;
      VIA 11.6 157.76 via_1600x480 ;
      VIA 334.8 152.32 via3_1600x480 ;
      VIA 334.8 152.32 via2_1600x480 ;
      VIA 334.8 152.32 via_1600x480 ;
      VIA 314.6 152.32 via3_1600x480 ;
      VIA 314.6 152.32 via2_1600x480 ;
      VIA 314.6 152.32 via_1600x480 ;
      VIA 294.4 152.32 via3_1600x480 ;
      VIA 294.4 152.32 via2_1600x480 ;
      VIA 294.4 152.32 via_1600x480 ;
      VIA 274.2 152.32 via3_1600x480 ;
      VIA 274.2 152.32 via2_1600x480 ;
      VIA 274.2 152.32 via_1600x480 ;
      VIA 254 152.32 via3_1600x480 ;
      VIA 254 152.32 via2_1600x480 ;
      VIA 254 152.32 via_1600x480 ;
      VIA 233.8 152.32 via3_1600x480 ;
      VIA 233.8 152.32 via2_1600x480 ;
      VIA 233.8 152.32 via_1600x480 ;
      VIA 213.6 152.32 via3_1600x480 ;
      VIA 213.6 152.32 via2_1600x480 ;
      VIA 213.6 152.32 via_1600x480 ;
      VIA 193.4 152.32 via3_1600x480 ;
      VIA 193.4 152.32 via2_1600x480 ;
      VIA 193.4 152.32 via_1600x480 ;
      VIA 173.2 152.32 via3_1600x480 ;
      VIA 173.2 152.32 via2_1600x480 ;
      VIA 173.2 152.32 via_1600x480 ;
      VIA 153 152.32 via3_1600x480 ;
      VIA 153 152.32 via2_1600x480 ;
      VIA 153 152.32 via_1600x480 ;
      VIA 132.8 152.32 via3_1600x480 ;
      VIA 132.8 152.32 via2_1600x480 ;
      VIA 132.8 152.32 via_1600x480 ;
      VIA 112.6 152.32 via3_1600x480 ;
      VIA 112.6 152.32 via2_1600x480 ;
      VIA 112.6 152.32 via_1600x480 ;
      VIA 92.4 152.32 via3_1600x480 ;
      VIA 92.4 152.32 via2_1600x480 ;
      VIA 92.4 152.32 via_1600x480 ;
      VIA 72.2 152.32 via3_1600x480 ;
      VIA 72.2 152.32 via2_1600x480 ;
      VIA 72.2 152.32 via_1600x480 ;
      VIA 52 152.32 via3_1600x480 ;
      VIA 52 152.32 via2_1600x480 ;
      VIA 52 152.32 via_1600x480 ;
      VIA 31.8 152.32 via3_1600x480 ;
      VIA 31.8 152.32 via2_1600x480 ;
      VIA 31.8 152.32 via_1600x480 ;
      VIA 11.6 152.32 via3_1600x480 ;
      VIA 11.6 152.32 via2_1600x480 ;
      VIA 11.6 152.32 via_1600x480 ;
      VIA 334.8 146.88 via3_1600x480 ;
      VIA 334.8 146.88 via2_1600x480 ;
      VIA 334.8 146.88 via_1600x480 ;
      VIA 314.6 146.88 via3_1600x480 ;
      VIA 314.6 146.88 via2_1600x480 ;
      VIA 314.6 146.88 via_1600x480 ;
      VIA 294.4 146.88 via3_1600x480 ;
      VIA 294.4 146.88 via2_1600x480 ;
      VIA 294.4 146.88 via_1600x480 ;
      VIA 274.2 146.88 via3_1600x480 ;
      VIA 274.2 146.88 via2_1600x480 ;
      VIA 274.2 146.88 via_1600x480 ;
      VIA 254 146.88 via3_1600x480 ;
      VIA 254 146.88 via2_1600x480 ;
      VIA 254 146.88 via_1600x480 ;
      VIA 233.8 146.88 via3_1600x480 ;
      VIA 233.8 146.88 via2_1600x480 ;
      VIA 233.8 146.88 via_1600x480 ;
      VIA 213.6 146.88 via3_1600x480 ;
      VIA 213.6 146.88 via2_1600x480 ;
      VIA 213.6 146.88 via_1600x480 ;
      VIA 193.4 146.88 via3_1600x480 ;
      VIA 193.4 146.88 via2_1600x480 ;
      VIA 193.4 146.88 via_1600x480 ;
      VIA 173.2 146.88 via3_1600x480 ;
      VIA 173.2 146.88 via2_1600x480 ;
      VIA 173.2 146.88 via_1600x480 ;
      VIA 153 146.88 via3_1600x480 ;
      VIA 153 146.88 via2_1600x480 ;
      VIA 153 146.88 via_1600x480 ;
      VIA 132.8 146.88 via3_1600x480 ;
      VIA 132.8 146.88 via2_1600x480 ;
      VIA 132.8 146.88 via_1600x480 ;
      VIA 112.6 146.88 via3_1600x480 ;
      VIA 112.6 146.88 via2_1600x480 ;
      VIA 112.6 146.88 via_1600x480 ;
      VIA 92.4 146.88 via3_1600x480 ;
      VIA 92.4 146.88 via2_1600x480 ;
      VIA 92.4 146.88 via_1600x480 ;
      VIA 72.2 146.88 via3_1600x480 ;
      VIA 72.2 146.88 via2_1600x480 ;
      VIA 72.2 146.88 via_1600x480 ;
      VIA 52 146.88 via3_1600x480 ;
      VIA 52 146.88 via2_1600x480 ;
      VIA 52 146.88 via_1600x480 ;
      VIA 31.8 146.88 via3_1600x480 ;
      VIA 31.8 146.88 via2_1600x480 ;
      VIA 31.8 146.88 via_1600x480 ;
      VIA 11.6 146.88 via3_1600x480 ;
      VIA 11.6 146.88 via2_1600x480 ;
      VIA 11.6 146.88 via_1600x480 ;
      VIA 334.8 141.44 via3_1600x480 ;
      VIA 334.8 141.44 via2_1600x480 ;
      VIA 334.8 141.44 via_1600x480 ;
      VIA 314.6 141.44 via3_1600x480 ;
      VIA 314.6 141.44 via2_1600x480 ;
      VIA 314.6 141.44 via_1600x480 ;
      VIA 294.4 141.44 via3_1600x480 ;
      VIA 294.4 141.44 via2_1600x480 ;
      VIA 294.4 141.44 via_1600x480 ;
      VIA 274.2 141.44 via3_1600x480 ;
      VIA 274.2 141.44 via2_1600x480 ;
      VIA 274.2 141.44 via_1600x480 ;
      VIA 254 141.44 via3_1600x480 ;
      VIA 254 141.44 via2_1600x480 ;
      VIA 254 141.44 via_1600x480 ;
      VIA 233.8 141.44 via3_1600x480 ;
      VIA 233.8 141.44 via2_1600x480 ;
      VIA 233.8 141.44 via_1600x480 ;
      VIA 213.6 141.44 via3_1600x480 ;
      VIA 213.6 141.44 via2_1600x480 ;
      VIA 213.6 141.44 via_1600x480 ;
      VIA 193.4 141.44 via3_1600x480 ;
      VIA 193.4 141.44 via2_1600x480 ;
      VIA 193.4 141.44 via_1600x480 ;
      VIA 173.2 141.44 via3_1600x480 ;
      VIA 173.2 141.44 via2_1600x480 ;
      VIA 173.2 141.44 via_1600x480 ;
      VIA 153 141.44 via3_1600x480 ;
      VIA 153 141.44 via2_1600x480 ;
      VIA 153 141.44 via_1600x480 ;
      VIA 132.8 141.44 via3_1600x480 ;
      VIA 132.8 141.44 via2_1600x480 ;
      VIA 132.8 141.44 via_1600x480 ;
      VIA 112.6 141.44 via3_1600x480 ;
      VIA 112.6 141.44 via2_1600x480 ;
      VIA 112.6 141.44 via_1600x480 ;
      VIA 92.4 141.44 via3_1600x480 ;
      VIA 92.4 141.44 via2_1600x480 ;
      VIA 92.4 141.44 via_1600x480 ;
      VIA 72.2 141.44 via3_1600x480 ;
      VIA 72.2 141.44 via2_1600x480 ;
      VIA 72.2 141.44 via_1600x480 ;
      VIA 52 141.44 via3_1600x480 ;
      VIA 52 141.44 via2_1600x480 ;
      VIA 52 141.44 via_1600x480 ;
      VIA 31.8 141.44 via3_1600x480 ;
      VIA 31.8 141.44 via2_1600x480 ;
      VIA 31.8 141.44 via_1600x480 ;
      VIA 11.6 141.44 via3_1600x480 ;
      VIA 11.6 141.44 via2_1600x480 ;
      VIA 11.6 141.44 via_1600x480 ;
      VIA 334.8 136 via3_1600x480 ;
      VIA 334.8 136 via2_1600x480 ;
      VIA 334.8 136 via_1600x480 ;
      VIA 314.6 136 via3_1600x480 ;
      VIA 314.6 136 via2_1600x480 ;
      VIA 314.6 136 via_1600x480 ;
      VIA 294.4 136 via3_1600x480 ;
      VIA 294.4 136 via2_1600x480 ;
      VIA 294.4 136 via_1600x480 ;
      VIA 274.2 136 via3_1600x480 ;
      VIA 274.2 136 via2_1600x480 ;
      VIA 274.2 136 via_1600x480 ;
      VIA 254 136 via3_1600x480 ;
      VIA 254 136 via2_1600x480 ;
      VIA 254 136 via_1600x480 ;
      VIA 233.8 136 via3_1600x480 ;
      VIA 233.8 136 via2_1600x480 ;
      VIA 233.8 136 via_1600x480 ;
      VIA 213.6 136 via3_1600x480 ;
      VIA 213.6 136 via2_1600x480 ;
      VIA 213.6 136 via_1600x480 ;
      VIA 193.4 136 via3_1600x480 ;
      VIA 193.4 136 via2_1600x480 ;
      VIA 193.4 136 via_1600x480 ;
      VIA 173.2 136 via3_1600x480 ;
      VIA 173.2 136 via2_1600x480 ;
      VIA 173.2 136 via_1600x480 ;
      VIA 153 136 via3_1600x480 ;
      VIA 153 136 via2_1600x480 ;
      VIA 153 136 via_1600x480 ;
      VIA 132.8 136 via3_1600x480 ;
      VIA 132.8 136 via2_1600x480 ;
      VIA 132.8 136 via_1600x480 ;
      VIA 112.6 136 via3_1600x480 ;
      VIA 112.6 136 via2_1600x480 ;
      VIA 112.6 136 via_1600x480 ;
      VIA 92.4 136 via3_1600x480 ;
      VIA 92.4 136 via2_1600x480 ;
      VIA 92.4 136 via_1600x480 ;
      VIA 72.2 136 via3_1600x480 ;
      VIA 72.2 136 via2_1600x480 ;
      VIA 72.2 136 via_1600x480 ;
      VIA 52 136 via3_1600x480 ;
      VIA 52 136 via2_1600x480 ;
      VIA 52 136 via_1600x480 ;
      VIA 31.8 136 via3_1600x480 ;
      VIA 31.8 136 via2_1600x480 ;
      VIA 31.8 136 via_1600x480 ;
      VIA 11.6 136 via3_1600x480 ;
      VIA 11.6 136 via2_1600x480 ;
      VIA 11.6 136 via_1600x480 ;
      VIA 334.8 130.56 via3_1600x480 ;
      VIA 334.8 130.56 via2_1600x480 ;
      VIA 334.8 130.56 via_1600x480 ;
      VIA 314.6 130.56 via3_1600x480 ;
      VIA 314.6 130.56 via2_1600x480 ;
      VIA 314.6 130.56 via_1600x480 ;
      VIA 294.4 130.56 via3_1600x480 ;
      VIA 294.4 130.56 via2_1600x480 ;
      VIA 294.4 130.56 via_1600x480 ;
      VIA 274.2 130.56 via3_1600x480 ;
      VIA 274.2 130.56 via2_1600x480 ;
      VIA 274.2 130.56 via_1600x480 ;
      VIA 254 130.56 via3_1600x480 ;
      VIA 254 130.56 via2_1600x480 ;
      VIA 254 130.56 via_1600x480 ;
      VIA 233.8 130.56 via3_1600x480 ;
      VIA 233.8 130.56 via2_1600x480 ;
      VIA 233.8 130.56 via_1600x480 ;
      VIA 213.6 130.56 via3_1600x480 ;
      VIA 213.6 130.56 via2_1600x480 ;
      VIA 213.6 130.56 via_1600x480 ;
      VIA 193.4 130.56 via3_1600x480 ;
      VIA 193.4 130.56 via2_1600x480 ;
      VIA 193.4 130.56 via_1600x480 ;
      VIA 173.2 130.56 via3_1600x480 ;
      VIA 173.2 130.56 via2_1600x480 ;
      VIA 173.2 130.56 via_1600x480 ;
      VIA 153 130.56 via3_1600x480 ;
      VIA 153 130.56 via2_1600x480 ;
      VIA 153 130.56 via_1600x480 ;
      VIA 132.8 130.56 via3_1600x480 ;
      VIA 132.8 130.56 via2_1600x480 ;
      VIA 132.8 130.56 via_1600x480 ;
      VIA 112.6 130.56 via3_1600x480 ;
      VIA 112.6 130.56 via2_1600x480 ;
      VIA 112.6 130.56 via_1600x480 ;
      VIA 92.4 130.56 via3_1600x480 ;
      VIA 92.4 130.56 via2_1600x480 ;
      VIA 92.4 130.56 via_1600x480 ;
      VIA 72.2 130.56 via3_1600x480 ;
      VIA 72.2 130.56 via2_1600x480 ;
      VIA 72.2 130.56 via_1600x480 ;
      VIA 52 130.56 via3_1600x480 ;
      VIA 52 130.56 via2_1600x480 ;
      VIA 52 130.56 via_1600x480 ;
      VIA 31.8 130.56 via3_1600x480 ;
      VIA 31.8 130.56 via2_1600x480 ;
      VIA 31.8 130.56 via_1600x480 ;
      VIA 11.6 130.56 via3_1600x480 ;
      VIA 11.6 130.56 via2_1600x480 ;
      VIA 11.6 130.56 via_1600x480 ;
      VIA 334.8 125.12 via3_1600x480 ;
      VIA 334.8 125.12 via2_1600x480 ;
      VIA 334.8 125.12 via_1600x480 ;
      VIA 314.6 125.12 via3_1600x480 ;
      VIA 314.6 125.12 via2_1600x480 ;
      VIA 314.6 125.12 via_1600x480 ;
      VIA 294.4 125.12 via3_1600x480 ;
      VIA 294.4 125.12 via2_1600x480 ;
      VIA 294.4 125.12 via_1600x480 ;
      VIA 274.2 125.12 via3_1600x480 ;
      VIA 274.2 125.12 via2_1600x480 ;
      VIA 274.2 125.12 via_1600x480 ;
      VIA 254 125.12 via3_1600x480 ;
      VIA 254 125.12 via2_1600x480 ;
      VIA 254 125.12 via_1600x480 ;
      VIA 233.8 125.12 via3_1600x480 ;
      VIA 233.8 125.12 via2_1600x480 ;
      VIA 233.8 125.12 via_1600x480 ;
      VIA 213.6 125.12 via3_1600x480 ;
      VIA 213.6 125.12 via2_1600x480 ;
      VIA 213.6 125.12 via_1600x480 ;
      VIA 193.4 125.12 via3_1600x480 ;
      VIA 193.4 125.12 via2_1600x480 ;
      VIA 193.4 125.12 via_1600x480 ;
      VIA 173.2 125.12 via3_1600x480 ;
      VIA 173.2 125.12 via2_1600x480 ;
      VIA 173.2 125.12 via_1600x480 ;
      VIA 153 125.12 via3_1600x480 ;
      VIA 153 125.12 via2_1600x480 ;
      VIA 153 125.12 via_1600x480 ;
      VIA 132.8 125.12 via3_1600x480 ;
      VIA 132.8 125.12 via2_1600x480 ;
      VIA 132.8 125.12 via_1600x480 ;
      VIA 112.6 125.12 via3_1600x480 ;
      VIA 112.6 125.12 via2_1600x480 ;
      VIA 112.6 125.12 via_1600x480 ;
      VIA 92.4 125.12 via3_1600x480 ;
      VIA 92.4 125.12 via2_1600x480 ;
      VIA 92.4 125.12 via_1600x480 ;
      VIA 72.2 125.12 via3_1600x480 ;
      VIA 72.2 125.12 via2_1600x480 ;
      VIA 72.2 125.12 via_1600x480 ;
      VIA 52 125.12 via3_1600x480 ;
      VIA 52 125.12 via2_1600x480 ;
      VIA 52 125.12 via_1600x480 ;
      VIA 31.8 125.12 via3_1600x480 ;
      VIA 31.8 125.12 via2_1600x480 ;
      VIA 31.8 125.12 via_1600x480 ;
      VIA 11.6 125.12 via3_1600x480 ;
      VIA 11.6 125.12 via2_1600x480 ;
      VIA 11.6 125.12 via_1600x480 ;
      VIA 334.8 119.68 via3_1600x480 ;
      VIA 334.8 119.68 via2_1600x480 ;
      VIA 334.8 119.68 via_1600x480 ;
      VIA 314.6 119.68 via3_1600x480 ;
      VIA 314.6 119.68 via2_1600x480 ;
      VIA 314.6 119.68 via_1600x480 ;
      VIA 294.4 119.68 via3_1600x480 ;
      VIA 294.4 119.68 via2_1600x480 ;
      VIA 294.4 119.68 via_1600x480 ;
      VIA 274.2 119.68 via3_1600x480 ;
      VIA 274.2 119.68 via2_1600x480 ;
      VIA 274.2 119.68 via_1600x480 ;
      VIA 254 119.68 via3_1600x480 ;
      VIA 254 119.68 via2_1600x480 ;
      VIA 254 119.68 via_1600x480 ;
      VIA 233.8 119.68 via3_1600x480 ;
      VIA 233.8 119.68 via2_1600x480 ;
      VIA 233.8 119.68 via_1600x480 ;
      VIA 213.6 119.68 via3_1600x480 ;
      VIA 213.6 119.68 via2_1600x480 ;
      VIA 213.6 119.68 via_1600x480 ;
      VIA 193.4 119.68 via3_1600x480 ;
      VIA 193.4 119.68 via2_1600x480 ;
      VIA 193.4 119.68 via_1600x480 ;
      VIA 173.2 119.68 via3_1600x480 ;
      VIA 173.2 119.68 via2_1600x480 ;
      VIA 173.2 119.68 via_1600x480 ;
      VIA 153 119.68 via3_1600x480 ;
      VIA 153 119.68 via2_1600x480 ;
      VIA 153 119.68 via_1600x480 ;
      VIA 132.8 119.68 via3_1600x480 ;
      VIA 132.8 119.68 via2_1600x480 ;
      VIA 132.8 119.68 via_1600x480 ;
      VIA 112.6 119.68 via3_1600x480 ;
      VIA 112.6 119.68 via2_1600x480 ;
      VIA 112.6 119.68 via_1600x480 ;
      VIA 92.4 119.68 via3_1600x480 ;
      VIA 92.4 119.68 via2_1600x480 ;
      VIA 92.4 119.68 via_1600x480 ;
      VIA 72.2 119.68 via3_1600x480 ;
      VIA 72.2 119.68 via2_1600x480 ;
      VIA 72.2 119.68 via_1600x480 ;
      VIA 52 119.68 via3_1600x480 ;
      VIA 52 119.68 via2_1600x480 ;
      VIA 52 119.68 via_1600x480 ;
      VIA 31.8 119.68 via3_1600x480 ;
      VIA 31.8 119.68 via2_1600x480 ;
      VIA 31.8 119.68 via_1600x480 ;
      VIA 11.6 119.68 via3_1600x480 ;
      VIA 11.6 119.68 via2_1600x480 ;
      VIA 11.6 119.68 via_1600x480 ;
      VIA 334.8 114.24 via3_1600x480 ;
      VIA 334.8 114.24 via2_1600x480 ;
      VIA 334.8 114.24 via_1600x480 ;
      VIA 314.6 114.24 via3_1600x480 ;
      VIA 314.6 114.24 via2_1600x480 ;
      VIA 314.6 114.24 via_1600x480 ;
      VIA 294.4 114.24 via3_1600x480 ;
      VIA 294.4 114.24 via2_1600x480 ;
      VIA 294.4 114.24 via_1600x480 ;
      VIA 274.2 114.24 via3_1600x480 ;
      VIA 274.2 114.24 via2_1600x480 ;
      VIA 274.2 114.24 via_1600x480 ;
      VIA 254 114.24 via3_1600x480 ;
      VIA 254 114.24 via2_1600x480 ;
      VIA 254 114.24 via_1600x480 ;
      VIA 233.8 114.24 via3_1600x480 ;
      VIA 233.8 114.24 via2_1600x480 ;
      VIA 233.8 114.24 via_1600x480 ;
      VIA 213.6 114.24 via3_1600x480 ;
      VIA 213.6 114.24 via2_1600x480 ;
      VIA 213.6 114.24 via_1600x480 ;
      VIA 193.4 114.24 via3_1600x480 ;
      VIA 193.4 114.24 via2_1600x480 ;
      VIA 193.4 114.24 via_1600x480 ;
      VIA 173.2 114.24 via3_1600x480 ;
      VIA 173.2 114.24 via2_1600x480 ;
      VIA 173.2 114.24 via_1600x480 ;
      VIA 153 114.24 via3_1600x480 ;
      VIA 153 114.24 via2_1600x480 ;
      VIA 153 114.24 via_1600x480 ;
      VIA 132.8 114.24 via3_1600x480 ;
      VIA 132.8 114.24 via2_1600x480 ;
      VIA 132.8 114.24 via_1600x480 ;
      VIA 112.6 114.24 via3_1600x480 ;
      VIA 112.6 114.24 via2_1600x480 ;
      VIA 112.6 114.24 via_1600x480 ;
      VIA 92.4 114.24 via3_1600x480 ;
      VIA 92.4 114.24 via2_1600x480 ;
      VIA 92.4 114.24 via_1600x480 ;
      VIA 72.2 114.24 via3_1600x480 ;
      VIA 72.2 114.24 via2_1600x480 ;
      VIA 72.2 114.24 via_1600x480 ;
      VIA 52 114.24 via3_1600x480 ;
      VIA 52 114.24 via2_1600x480 ;
      VIA 52 114.24 via_1600x480 ;
      VIA 31.8 114.24 via3_1600x480 ;
      VIA 31.8 114.24 via2_1600x480 ;
      VIA 31.8 114.24 via_1600x480 ;
      VIA 11.6 114.24 via3_1600x480 ;
      VIA 11.6 114.24 via2_1600x480 ;
      VIA 11.6 114.24 via_1600x480 ;
      VIA 334.8 108.8 via3_1600x480 ;
      VIA 334.8 108.8 via2_1600x480 ;
      VIA 334.8 108.8 via_1600x480 ;
      VIA 314.6 108.8 via3_1600x480 ;
      VIA 314.6 108.8 via2_1600x480 ;
      VIA 314.6 108.8 via_1600x480 ;
      VIA 294.4 108.8 via3_1600x480 ;
      VIA 294.4 108.8 via2_1600x480 ;
      VIA 294.4 108.8 via_1600x480 ;
      VIA 274.2 108.8 via3_1600x480 ;
      VIA 274.2 108.8 via2_1600x480 ;
      VIA 274.2 108.8 via_1600x480 ;
      VIA 254 108.8 via3_1600x480 ;
      VIA 254 108.8 via2_1600x480 ;
      VIA 254 108.8 via_1600x480 ;
      VIA 233.8 108.8 via3_1600x480 ;
      VIA 233.8 108.8 via2_1600x480 ;
      VIA 233.8 108.8 via_1600x480 ;
      VIA 213.6 108.8 via3_1600x480 ;
      VIA 213.6 108.8 via2_1600x480 ;
      VIA 213.6 108.8 via_1600x480 ;
      VIA 193.4 108.8 via3_1600x480 ;
      VIA 193.4 108.8 via2_1600x480 ;
      VIA 193.4 108.8 via_1600x480 ;
      VIA 173.2 108.8 via3_1600x480 ;
      VIA 173.2 108.8 via2_1600x480 ;
      VIA 173.2 108.8 via_1600x480 ;
      VIA 153 108.8 via3_1600x480 ;
      VIA 153 108.8 via2_1600x480 ;
      VIA 153 108.8 via_1600x480 ;
      VIA 132.8 108.8 via3_1600x480 ;
      VIA 132.8 108.8 via2_1600x480 ;
      VIA 132.8 108.8 via_1600x480 ;
      VIA 112.6 108.8 via3_1600x480 ;
      VIA 112.6 108.8 via2_1600x480 ;
      VIA 112.6 108.8 via_1600x480 ;
      VIA 92.4 108.8 via3_1600x480 ;
      VIA 92.4 108.8 via2_1600x480 ;
      VIA 92.4 108.8 via_1600x480 ;
      VIA 72.2 108.8 via3_1600x480 ;
      VIA 72.2 108.8 via2_1600x480 ;
      VIA 72.2 108.8 via_1600x480 ;
      VIA 52 108.8 via3_1600x480 ;
      VIA 52 108.8 via2_1600x480 ;
      VIA 52 108.8 via_1600x480 ;
      VIA 31.8 108.8 via3_1600x480 ;
      VIA 31.8 108.8 via2_1600x480 ;
      VIA 31.8 108.8 via_1600x480 ;
      VIA 11.6 108.8 via3_1600x480 ;
      VIA 11.6 108.8 via2_1600x480 ;
      VIA 11.6 108.8 via_1600x480 ;
      VIA 334.8 103.36 via3_1600x480 ;
      VIA 334.8 103.36 via2_1600x480 ;
      VIA 334.8 103.36 via_1600x480 ;
      VIA 314.6 103.36 via3_1600x480 ;
      VIA 314.6 103.36 via2_1600x480 ;
      VIA 314.6 103.36 via_1600x480 ;
      VIA 294.4 103.36 via3_1600x480 ;
      VIA 294.4 103.36 via2_1600x480 ;
      VIA 294.4 103.36 via_1600x480 ;
      VIA 274.2 103.36 via3_1600x480 ;
      VIA 274.2 103.36 via2_1600x480 ;
      VIA 274.2 103.36 via_1600x480 ;
      VIA 254 103.36 via3_1600x480 ;
      VIA 254 103.36 via2_1600x480 ;
      VIA 254 103.36 via_1600x480 ;
      VIA 233.8 103.36 via3_1600x480 ;
      VIA 233.8 103.36 via2_1600x480 ;
      VIA 233.8 103.36 via_1600x480 ;
      VIA 213.6 103.36 via3_1600x480 ;
      VIA 213.6 103.36 via2_1600x480 ;
      VIA 213.6 103.36 via_1600x480 ;
      VIA 193.4 103.36 via3_1600x480 ;
      VIA 193.4 103.36 via2_1600x480 ;
      VIA 193.4 103.36 via_1600x480 ;
      VIA 173.2 103.36 via3_1600x480 ;
      VIA 173.2 103.36 via2_1600x480 ;
      VIA 173.2 103.36 via_1600x480 ;
      VIA 153 103.36 via3_1600x480 ;
      VIA 153 103.36 via2_1600x480 ;
      VIA 153 103.36 via_1600x480 ;
      VIA 132.8 103.36 via3_1600x480 ;
      VIA 132.8 103.36 via2_1600x480 ;
      VIA 132.8 103.36 via_1600x480 ;
      VIA 112.6 103.36 via3_1600x480 ;
      VIA 112.6 103.36 via2_1600x480 ;
      VIA 112.6 103.36 via_1600x480 ;
      VIA 92.4 103.36 via3_1600x480 ;
      VIA 92.4 103.36 via2_1600x480 ;
      VIA 92.4 103.36 via_1600x480 ;
      VIA 72.2 103.36 via3_1600x480 ;
      VIA 72.2 103.36 via2_1600x480 ;
      VIA 72.2 103.36 via_1600x480 ;
      VIA 52 103.36 via3_1600x480 ;
      VIA 52 103.36 via2_1600x480 ;
      VIA 52 103.36 via_1600x480 ;
      VIA 31.8 103.36 via3_1600x480 ;
      VIA 31.8 103.36 via2_1600x480 ;
      VIA 31.8 103.36 via_1600x480 ;
      VIA 11.6 103.36 via3_1600x480 ;
      VIA 11.6 103.36 via2_1600x480 ;
      VIA 11.6 103.36 via_1600x480 ;
      VIA 334.8 97.92 via3_1600x480 ;
      VIA 334.8 97.92 via2_1600x480 ;
      VIA 334.8 97.92 via_1600x480 ;
      VIA 314.6 97.92 via3_1600x480 ;
      VIA 314.6 97.92 via2_1600x480 ;
      VIA 314.6 97.92 via_1600x480 ;
      VIA 294.4 97.92 via3_1600x480 ;
      VIA 294.4 97.92 via2_1600x480 ;
      VIA 294.4 97.92 via_1600x480 ;
      VIA 274.2 97.92 via3_1600x480 ;
      VIA 274.2 97.92 via2_1600x480 ;
      VIA 274.2 97.92 via_1600x480 ;
      VIA 254 97.92 via3_1600x480 ;
      VIA 254 97.92 via2_1600x480 ;
      VIA 254 97.92 via_1600x480 ;
      VIA 233.8 97.92 via3_1600x480 ;
      VIA 233.8 97.92 via2_1600x480 ;
      VIA 233.8 97.92 via_1600x480 ;
      VIA 213.6 97.92 via3_1600x480 ;
      VIA 213.6 97.92 via2_1600x480 ;
      VIA 213.6 97.92 via_1600x480 ;
      VIA 193.4 97.92 via3_1600x480 ;
      VIA 193.4 97.92 via2_1600x480 ;
      VIA 193.4 97.92 via_1600x480 ;
      VIA 173.2 97.92 via3_1600x480 ;
      VIA 173.2 97.92 via2_1600x480 ;
      VIA 173.2 97.92 via_1600x480 ;
      VIA 153 97.92 via3_1600x480 ;
      VIA 153 97.92 via2_1600x480 ;
      VIA 153 97.92 via_1600x480 ;
      VIA 132.8 97.92 via3_1600x480 ;
      VIA 132.8 97.92 via2_1600x480 ;
      VIA 132.8 97.92 via_1600x480 ;
      VIA 112.6 97.92 via3_1600x480 ;
      VIA 112.6 97.92 via2_1600x480 ;
      VIA 112.6 97.92 via_1600x480 ;
      VIA 92.4 97.92 via3_1600x480 ;
      VIA 92.4 97.92 via2_1600x480 ;
      VIA 92.4 97.92 via_1600x480 ;
      VIA 72.2 97.92 via3_1600x480 ;
      VIA 72.2 97.92 via2_1600x480 ;
      VIA 72.2 97.92 via_1600x480 ;
      VIA 52 97.92 via3_1600x480 ;
      VIA 52 97.92 via2_1600x480 ;
      VIA 52 97.92 via_1600x480 ;
      VIA 31.8 97.92 via3_1600x480 ;
      VIA 31.8 97.92 via2_1600x480 ;
      VIA 31.8 97.92 via_1600x480 ;
      VIA 11.6 97.92 via3_1600x480 ;
      VIA 11.6 97.92 via2_1600x480 ;
      VIA 11.6 97.92 via_1600x480 ;
      VIA 334.8 92.48 via3_1600x480 ;
      VIA 334.8 92.48 via2_1600x480 ;
      VIA 334.8 92.48 via_1600x480 ;
      VIA 314.6 92.48 via3_1600x480 ;
      VIA 314.6 92.48 via2_1600x480 ;
      VIA 314.6 92.48 via_1600x480 ;
      VIA 294.4 92.48 via3_1600x480 ;
      VIA 294.4 92.48 via2_1600x480 ;
      VIA 294.4 92.48 via_1600x480 ;
      VIA 274.2 92.48 via3_1600x480 ;
      VIA 274.2 92.48 via2_1600x480 ;
      VIA 274.2 92.48 via_1600x480 ;
      VIA 254 92.48 via3_1600x480 ;
      VIA 254 92.48 via2_1600x480 ;
      VIA 254 92.48 via_1600x480 ;
      VIA 233.8 92.48 via3_1600x480 ;
      VIA 233.8 92.48 via2_1600x480 ;
      VIA 233.8 92.48 via_1600x480 ;
      VIA 213.6 92.48 via3_1600x480 ;
      VIA 213.6 92.48 via2_1600x480 ;
      VIA 213.6 92.48 via_1600x480 ;
      VIA 193.4 92.48 via3_1600x480 ;
      VIA 193.4 92.48 via2_1600x480 ;
      VIA 193.4 92.48 via_1600x480 ;
      VIA 173.2 92.48 via3_1600x480 ;
      VIA 173.2 92.48 via2_1600x480 ;
      VIA 173.2 92.48 via_1600x480 ;
      VIA 153 92.48 via3_1600x480 ;
      VIA 153 92.48 via2_1600x480 ;
      VIA 153 92.48 via_1600x480 ;
      VIA 132.8 92.48 via3_1600x480 ;
      VIA 132.8 92.48 via2_1600x480 ;
      VIA 132.8 92.48 via_1600x480 ;
      VIA 112.6 92.48 via3_1600x480 ;
      VIA 112.6 92.48 via2_1600x480 ;
      VIA 112.6 92.48 via_1600x480 ;
      VIA 92.4 92.48 via3_1600x480 ;
      VIA 92.4 92.48 via2_1600x480 ;
      VIA 92.4 92.48 via_1600x480 ;
      VIA 72.2 92.48 via3_1600x480 ;
      VIA 72.2 92.48 via2_1600x480 ;
      VIA 72.2 92.48 via_1600x480 ;
      VIA 52 92.48 via3_1600x480 ;
      VIA 52 92.48 via2_1600x480 ;
      VIA 52 92.48 via_1600x480 ;
      VIA 31.8 92.48 via3_1600x480 ;
      VIA 31.8 92.48 via2_1600x480 ;
      VIA 31.8 92.48 via_1600x480 ;
      VIA 11.6 92.48 via3_1600x480 ;
      VIA 11.6 92.48 via2_1600x480 ;
      VIA 11.6 92.48 via_1600x480 ;
      VIA 334.8 87.04 via3_1600x480 ;
      VIA 334.8 87.04 via2_1600x480 ;
      VIA 334.8 87.04 via_1600x480 ;
      VIA 314.6 87.04 via3_1600x480 ;
      VIA 314.6 87.04 via2_1600x480 ;
      VIA 314.6 87.04 via_1600x480 ;
      VIA 294.4 87.04 via3_1600x480 ;
      VIA 294.4 87.04 via2_1600x480 ;
      VIA 294.4 87.04 via_1600x480 ;
      VIA 274.2 87.04 via3_1600x480 ;
      VIA 274.2 87.04 via2_1600x480 ;
      VIA 274.2 87.04 via_1600x480 ;
      VIA 254 87.04 via3_1600x480 ;
      VIA 254 87.04 via2_1600x480 ;
      VIA 254 87.04 via_1600x480 ;
      VIA 233.8 87.04 via3_1600x480 ;
      VIA 233.8 87.04 via2_1600x480 ;
      VIA 233.8 87.04 via_1600x480 ;
      VIA 213.6 87.04 via3_1600x480 ;
      VIA 213.6 87.04 via2_1600x480 ;
      VIA 213.6 87.04 via_1600x480 ;
      VIA 193.4 87.04 via3_1600x480 ;
      VIA 193.4 87.04 via2_1600x480 ;
      VIA 193.4 87.04 via_1600x480 ;
      VIA 173.2 87.04 via3_1600x480 ;
      VIA 173.2 87.04 via2_1600x480 ;
      VIA 173.2 87.04 via_1600x480 ;
      VIA 153 87.04 via3_1600x480 ;
      VIA 153 87.04 via2_1600x480 ;
      VIA 153 87.04 via_1600x480 ;
      VIA 132.8 87.04 via3_1600x480 ;
      VIA 132.8 87.04 via2_1600x480 ;
      VIA 132.8 87.04 via_1600x480 ;
      VIA 112.6 87.04 via3_1600x480 ;
      VIA 112.6 87.04 via2_1600x480 ;
      VIA 112.6 87.04 via_1600x480 ;
      VIA 92.4 87.04 via3_1600x480 ;
      VIA 92.4 87.04 via2_1600x480 ;
      VIA 92.4 87.04 via_1600x480 ;
      VIA 72.2 87.04 via3_1600x480 ;
      VIA 72.2 87.04 via2_1600x480 ;
      VIA 72.2 87.04 via_1600x480 ;
      VIA 52 87.04 via3_1600x480 ;
      VIA 52 87.04 via2_1600x480 ;
      VIA 52 87.04 via_1600x480 ;
      VIA 31.8 87.04 via3_1600x480 ;
      VIA 31.8 87.04 via2_1600x480 ;
      VIA 31.8 87.04 via_1600x480 ;
      VIA 11.6 87.04 via3_1600x480 ;
      VIA 11.6 87.04 via2_1600x480 ;
      VIA 11.6 87.04 via_1600x480 ;
      VIA 334.8 81.6 via3_1600x480 ;
      VIA 334.8 81.6 via2_1600x480 ;
      VIA 334.8 81.6 via_1600x480 ;
      VIA 314.6 81.6 via3_1600x480 ;
      VIA 314.6 81.6 via2_1600x480 ;
      VIA 314.6 81.6 via_1600x480 ;
      VIA 294.4 81.6 via3_1600x480 ;
      VIA 294.4 81.6 via2_1600x480 ;
      VIA 294.4 81.6 via_1600x480 ;
      VIA 274.2 81.6 via3_1600x480 ;
      VIA 274.2 81.6 via2_1600x480 ;
      VIA 274.2 81.6 via_1600x480 ;
      VIA 254 81.6 via3_1600x480 ;
      VIA 254 81.6 via2_1600x480 ;
      VIA 254 81.6 via_1600x480 ;
      VIA 233.8 81.6 via3_1600x480 ;
      VIA 233.8 81.6 via2_1600x480 ;
      VIA 233.8 81.6 via_1600x480 ;
      VIA 213.6 81.6 via3_1600x480 ;
      VIA 213.6 81.6 via2_1600x480 ;
      VIA 213.6 81.6 via_1600x480 ;
      VIA 193.4 81.6 via3_1600x480 ;
      VIA 193.4 81.6 via2_1600x480 ;
      VIA 193.4 81.6 via_1600x480 ;
      VIA 173.2 81.6 via3_1600x480 ;
      VIA 173.2 81.6 via2_1600x480 ;
      VIA 173.2 81.6 via_1600x480 ;
      VIA 153 81.6 via3_1600x480 ;
      VIA 153 81.6 via2_1600x480 ;
      VIA 153 81.6 via_1600x480 ;
      VIA 132.8 81.6 via3_1600x480 ;
      VIA 132.8 81.6 via2_1600x480 ;
      VIA 132.8 81.6 via_1600x480 ;
      VIA 112.6 81.6 via3_1600x480 ;
      VIA 112.6 81.6 via2_1600x480 ;
      VIA 112.6 81.6 via_1600x480 ;
      VIA 92.4 81.6 via3_1600x480 ;
      VIA 92.4 81.6 via2_1600x480 ;
      VIA 92.4 81.6 via_1600x480 ;
      VIA 72.2 81.6 via3_1600x480 ;
      VIA 72.2 81.6 via2_1600x480 ;
      VIA 72.2 81.6 via_1600x480 ;
      VIA 52 81.6 via3_1600x480 ;
      VIA 52 81.6 via2_1600x480 ;
      VIA 52 81.6 via_1600x480 ;
      VIA 31.8 81.6 via3_1600x480 ;
      VIA 31.8 81.6 via2_1600x480 ;
      VIA 31.8 81.6 via_1600x480 ;
      VIA 11.6 81.6 via3_1600x480 ;
      VIA 11.6 81.6 via2_1600x480 ;
      VIA 11.6 81.6 via_1600x480 ;
      VIA 334.8 76.16 via3_1600x480 ;
      VIA 334.8 76.16 via2_1600x480 ;
      VIA 334.8 76.16 via_1600x480 ;
      VIA 314.6 76.16 via3_1600x480 ;
      VIA 314.6 76.16 via2_1600x480 ;
      VIA 314.6 76.16 via_1600x480 ;
      VIA 294.4 76.16 via3_1600x480 ;
      VIA 294.4 76.16 via2_1600x480 ;
      VIA 294.4 76.16 via_1600x480 ;
      VIA 274.2 76.16 via3_1600x480 ;
      VIA 274.2 76.16 via2_1600x480 ;
      VIA 274.2 76.16 via_1600x480 ;
      VIA 254 76.16 via3_1600x480 ;
      VIA 254 76.16 via2_1600x480 ;
      VIA 254 76.16 via_1600x480 ;
      VIA 233.8 76.16 via3_1600x480 ;
      VIA 233.8 76.16 via2_1600x480 ;
      VIA 233.8 76.16 via_1600x480 ;
      VIA 213.6 76.16 via3_1600x480 ;
      VIA 213.6 76.16 via2_1600x480 ;
      VIA 213.6 76.16 via_1600x480 ;
      VIA 193.4 76.16 via3_1600x480 ;
      VIA 193.4 76.16 via2_1600x480 ;
      VIA 193.4 76.16 via_1600x480 ;
      VIA 173.2 76.16 via3_1600x480 ;
      VIA 173.2 76.16 via2_1600x480 ;
      VIA 173.2 76.16 via_1600x480 ;
      VIA 153 76.16 via3_1600x480 ;
      VIA 153 76.16 via2_1600x480 ;
      VIA 153 76.16 via_1600x480 ;
      VIA 132.8 76.16 via3_1600x480 ;
      VIA 132.8 76.16 via2_1600x480 ;
      VIA 132.8 76.16 via_1600x480 ;
      VIA 112.6 76.16 via3_1600x480 ;
      VIA 112.6 76.16 via2_1600x480 ;
      VIA 112.6 76.16 via_1600x480 ;
      VIA 92.4 76.16 via3_1600x480 ;
      VIA 92.4 76.16 via2_1600x480 ;
      VIA 92.4 76.16 via_1600x480 ;
      VIA 72.2 76.16 via3_1600x480 ;
      VIA 72.2 76.16 via2_1600x480 ;
      VIA 72.2 76.16 via_1600x480 ;
      VIA 52 76.16 via3_1600x480 ;
      VIA 52 76.16 via2_1600x480 ;
      VIA 52 76.16 via_1600x480 ;
      VIA 31.8 76.16 via3_1600x480 ;
      VIA 31.8 76.16 via2_1600x480 ;
      VIA 31.8 76.16 via_1600x480 ;
      VIA 11.6 76.16 via3_1600x480 ;
      VIA 11.6 76.16 via2_1600x480 ;
      VIA 11.6 76.16 via_1600x480 ;
      VIA 334.8 70.72 via3_1600x480 ;
      VIA 334.8 70.72 via2_1600x480 ;
      VIA 334.8 70.72 via_1600x480 ;
      VIA 314.6 70.72 via3_1600x480 ;
      VIA 314.6 70.72 via2_1600x480 ;
      VIA 314.6 70.72 via_1600x480 ;
      VIA 294.4 70.72 via3_1600x480 ;
      VIA 294.4 70.72 via2_1600x480 ;
      VIA 294.4 70.72 via_1600x480 ;
      VIA 274.2 70.72 via3_1600x480 ;
      VIA 274.2 70.72 via2_1600x480 ;
      VIA 274.2 70.72 via_1600x480 ;
      VIA 254 70.72 via3_1600x480 ;
      VIA 254 70.72 via2_1600x480 ;
      VIA 254 70.72 via_1600x480 ;
      VIA 233.8 70.72 via3_1600x480 ;
      VIA 233.8 70.72 via2_1600x480 ;
      VIA 233.8 70.72 via_1600x480 ;
      VIA 213.6 70.72 via3_1600x480 ;
      VIA 213.6 70.72 via2_1600x480 ;
      VIA 213.6 70.72 via_1600x480 ;
      VIA 193.4 70.72 via3_1600x480 ;
      VIA 193.4 70.72 via2_1600x480 ;
      VIA 193.4 70.72 via_1600x480 ;
      VIA 173.2 70.72 via3_1600x480 ;
      VIA 173.2 70.72 via2_1600x480 ;
      VIA 173.2 70.72 via_1600x480 ;
      VIA 153 70.72 via3_1600x480 ;
      VIA 153 70.72 via2_1600x480 ;
      VIA 153 70.72 via_1600x480 ;
      VIA 132.8 70.72 via3_1600x480 ;
      VIA 132.8 70.72 via2_1600x480 ;
      VIA 132.8 70.72 via_1600x480 ;
      VIA 112.6 70.72 via3_1600x480 ;
      VIA 112.6 70.72 via2_1600x480 ;
      VIA 112.6 70.72 via_1600x480 ;
      VIA 92.4 70.72 via3_1600x480 ;
      VIA 92.4 70.72 via2_1600x480 ;
      VIA 92.4 70.72 via_1600x480 ;
      VIA 72.2 70.72 via3_1600x480 ;
      VIA 72.2 70.72 via2_1600x480 ;
      VIA 72.2 70.72 via_1600x480 ;
      VIA 52 70.72 via3_1600x480 ;
      VIA 52 70.72 via2_1600x480 ;
      VIA 52 70.72 via_1600x480 ;
      VIA 31.8 70.72 via3_1600x480 ;
      VIA 31.8 70.72 via2_1600x480 ;
      VIA 31.8 70.72 via_1600x480 ;
      VIA 11.6 70.72 via3_1600x480 ;
      VIA 11.6 70.72 via2_1600x480 ;
      VIA 11.6 70.72 via_1600x480 ;
      VIA 334.8 65.28 via3_1600x480 ;
      VIA 334.8 65.28 via2_1600x480 ;
      VIA 334.8 65.28 via_1600x480 ;
      VIA 314.6 65.28 via3_1600x480 ;
      VIA 314.6 65.28 via2_1600x480 ;
      VIA 314.6 65.28 via_1600x480 ;
      VIA 294.4 65.28 via3_1600x480 ;
      VIA 294.4 65.28 via2_1600x480 ;
      VIA 294.4 65.28 via_1600x480 ;
      VIA 274.2 65.28 via3_1600x480 ;
      VIA 274.2 65.28 via2_1600x480 ;
      VIA 274.2 65.28 via_1600x480 ;
      VIA 254 65.28 via3_1600x480 ;
      VIA 254 65.28 via2_1600x480 ;
      VIA 254 65.28 via_1600x480 ;
      VIA 233.8 65.28 via3_1600x480 ;
      VIA 233.8 65.28 via2_1600x480 ;
      VIA 233.8 65.28 via_1600x480 ;
      VIA 213.6 65.28 via3_1600x480 ;
      VIA 213.6 65.28 via2_1600x480 ;
      VIA 213.6 65.28 via_1600x480 ;
      VIA 193.4 65.28 via3_1600x480 ;
      VIA 193.4 65.28 via2_1600x480 ;
      VIA 193.4 65.28 via_1600x480 ;
      VIA 173.2 65.28 via3_1600x480 ;
      VIA 173.2 65.28 via2_1600x480 ;
      VIA 173.2 65.28 via_1600x480 ;
      VIA 153 65.28 via3_1600x480 ;
      VIA 153 65.28 via2_1600x480 ;
      VIA 153 65.28 via_1600x480 ;
      VIA 132.8 65.28 via3_1600x480 ;
      VIA 132.8 65.28 via2_1600x480 ;
      VIA 132.8 65.28 via_1600x480 ;
      VIA 112.6 65.28 via3_1600x480 ;
      VIA 112.6 65.28 via2_1600x480 ;
      VIA 112.6 65.28 via_1600x480 ;
      VIA 92.4 65.28 via3_1600x480 ;
      VIA 92.4 65.28 via2_1600x480 ;
      VIA 92.4 65.28 via_1600x480 ;
      VIA 72.2 65.28 via3_1600x480 ;
      VIA 72.2 65.28 via2_1600x480 ;
      VIA 72.2 65.28 via_1600x480 ;
      VIA 52 65.28 via3_1600x480 ;
      VIA 52 65.28 via2_1600x480 ;
      VIA 52 65.28 via_1600x480 ;
      VIA 31.8 65.28 via3_1600x480 ;
      VIA 31.8 65.28 via2_1600x480 ;
      VIA 31.8 65.28 via_1600x480 ;
      VIA 11.6 65.28 via3_1600x480 ;
      VIA 11.6 65.28 via2_1600x480 ;
      VIA 11.6 65.28 via_1600x480 ;
      VIA 334.8 59.84 via3_1600x480 ;
      VIA 334.8 59.84 via2_1600x480 ;
      VIA 334.8 59.84 via_1600x480 ;
      VIA 314.6 59.84 via3_1600x480 ;
      VIA 314.6 59.84 via2_1600x480 ;
      VIA 314.6 59.84 via_1600x480 ;
      VIA 294.4 59.84 via3_1600x480 ;
      VIA 294.4 59.84 via2_1600x480 ;
      VIA 294.4 59.84 via_1600x480 ;
      VIA 274.2 59.84 via3_1600x480 ;
      VIA 274.2 59.84 via2_1600x480 ;
      VIA 274.2 59.84 via_1600x480 ;
      VIA 254 59.84 via3_1600x480 ;
      VIA 254 59.84 via2_1600x480 ;
      VIA 254 59.84 via_1600x480 ;
      VIA 233.8 59.84 via3_1600x480 ;
      VIA 233.8 59.84 via2_1600x480 ;
      VIA 233.8 59.84 via_1600x480 ;
      VIA 213.6 59.84 via3_1600x480 ;
      VIA 213.6 59.84 via2_1600x480 ;
      VIA 213.6 59.84 via_1600x480 ;
      VIA 193.4 59.84 via3_1600x480 ;
      VIA 193.4 59.84 via2_1600x480 ;
      VIA 193.4 59.84 via_1600x480 ;
      VIA 173.2 59.84 via3_1600x480 ;
      VIA 173.2 59.84 via2_1600x480 ;
      VIA 173.2 59.84 via_1600x480 ;
      VIA 153 59.84 via3_1600x480 ;
      VIA 153 59.84 via2_1600x480 ;
      VIA 153 59.84 via_1600x480 ;
      VIA 132.8 59.84 via3_1600x480 ;
      VIA 132.8 59.84 via2_1600x480 ;
      VIA 132.8 59.84 via_1600x480 ;
      VIA 112.6 59.84 via3_1600x480 ;
      VIA 112.6 59.84 via2_1600x480 ;
      VIA 112.6 59.84 via_1600x480 ;
      VIA 92.4 59.84 via3_1600x480 ;
      VIA 92.4 59.84 via2_1600x480 ;
      VIA 92.4 59.84 via_1600x480 ;
      VIA 72.2 59.84 via3_1600x480 ;
      VIA 72.2 59.84 via2_1600x480 ;
      VIA 72.2 59.84 via_1600x480 ;
      VIA 52 59.84 via3_1600x480 ;
      VIA 52 59.84 via2_1600x480 ;
      VIA 52 59.84 via_1600x480 ;
      VIA 31.8 59.84 via3_1600x480 ;
      VIA 31.8 59.84 via2_1600x480 ;
      VIA 31.8 59.84 via_1600x480 ;
      VIA 11.6 59.84 via3_1600x480 ;
      VIA 11.6 59.84 via2_1600x480 ;
      VIA 11.6 59.84 via_1600x480 ;
      VIA 334.8 54.4 via3_1600x480 ;
      VIA 334.8 54.4 via2_1600x480 ;
      VIA 334.8 54.4 via_1600x480 ;
      VIA 314.6 54.4 via3_1600x480 ;
      VIA 314.6 54.4 via2_1600x480 ;
      VIA 314.6 54.4 via_1600x480 ;
      VIA 294.4 54.4 via3_1600x480 ;
      VIA 294.4 54.4 via2_1600x480 ;
      VIA 294.4 54.4 via_1600x480 ;
      VIA 274.2 54.4 via3_1600x480 ;
      VIA 274.2 54.4 via2_1600x480 ;
      VIA 274.2 54.4 via_1600x480 ;
      VIA 254 54.4 via3_1600x480 ;
      VIA 254 54.4 via2_1600x480 ;
      VIA 254 54.4 via_1600x480 ;
      VIA 233.8 54.4 via3_1600x480 ;
      VIA 233.8 54.4 via2_1600x480 ;
      VIA 233.8 54.4 via_1600x480 ;
      VIA 213.6 54.4 via3_1600x480 ;
      VIA 213.6 54.4 via2_1600x480 ;
      VIA 213.6 54.4 via_1600x480 ;
      VIA 193.4 54.4 via3_1600x480 ;
      VIA 193.4 54.4 via2_1600x480 ;
      VIA 193.4 54.4 via_1600x480 ;
      VIA 173.2 54.4 via3_1600x480 ;
      VIA 173.2 54.4 via2_1600x480 ;
      VIA 173.2 54.4 via_1600x480 ;
      VIA 153 54.4 via3_1600x480 ;
      VIA 153 54.4 via2_1600x480 ;
      VIA 153 54.4 via_1600x480 ;
      VIA 132.8 54.4 via3_1600x480 ;
      VIA 132.8 54.4 via2_1600x480 ;
      VIA 132.8 54.4 via_1600x480 ;
      VIA 112.6 54.4 via3_1600x480 ;
      VIA 112.6 54.4 via2_1600x480 ;
      VIA 112.6 54.4 via_1600x480 ;
      VIA 92.4 54.4 via3_1600x480 ;
      VIA 92.4 54.4 via2_1600x480 ;
      VIA 92.4 54.4 via_1600x480 ;
      VIA 72.2 54.4 via3_1600x480 ;
      VIA 72.2 54.4 via2_1600x480 ;
      VIA 72.2 54.4 via_1600x480 ;
      VIA 52 54.4 via3_1600x480 ;
      VIA 52 54.4 via2_1600x480 ;
      VIA 52 54.4 via_1600x480 ;
      VIA 31.8 54.4 via3_1600x480 ;
      VIA 31.8 54.4 via2_1600x480 ;
      VIA 31.8 54.4 via_1600x480 ;
      VIA 11.6 54.4 via3_1600x480 ;
      VIA 11.6 54.4 via2_1600x480 ;
      VIA 11.6 54.4 via_1600x480 ;
      VIA 334.8 48.96 via3_1600x480 ;
      VIA 334.8 48.96 via2_1600x480 ;
      VIA 334.8 48.96 via_1600x480 ;
      VIA 314.6 48.96 via3_1600x480 ;
      VIA 314.6 48.96 via2_1600x480 ;
      VIA 314.6 48.96 via_1600x480 ;
      VIA 294.4 48.96 via3_1600x480 ;
      VIA 294.4 48.96 via2_1600x480 ;
      VIA 294.4 48.96 via_1600x480 ;
      VIA 274.2 48.96 via3_1600x480 ;
      VIA 274.2 48.96 via2_1600x480 ;
      VIA 274.2 48.96 via_1600x480 ;
      VIA 254 48.96 via3_1600x480 ;
      VIA 254 48.96 via2_1600x480 ;
      VIA 254 48.96 via_1600x480 ;
      VIA 233.8 48.96 via3_1600x480 ;
      VIA 233.8 48.96 via2_1600x480 ;
      VIA 233.8 48.96 via_1600x480 ;
      VIA 213.6 48.96 via3_1600x480 ;
      VIA 213.6 48.96 via2_1600x480 ;
      VIA 213.6 48.96 via_1600x480 ;
      VIA 193.4 48.96 via3_1600x480 ;
      VIA 193.4 48.96 via2_1600x480 ;
      VIA 193.4 48.96 via_1600x480 ;
      VIA 173.2 48.96 via3_1600x480 ;
      VIA 173.2 48.96 via2_1600x480 ;
      VIA 173.2 48.96 via_1600x480 ;
      VIA 153 48.96 via3_1600x480 ;
      VIA 153 48.96 via2_1600x480 ;
      VIA 153 48.96 via_1600x480 ;
      VIA 132.8 48.96 via3_1600x480 ;
      VIA 132.8 48.96 via2_1600x480 ;
      VIA 132.8 48.96 via_1600x480 ;
      VIA 112.6 48.96 via3_1600x480 ;
      VIA 112.6 48.96 via2_1600x480 ;
      VIA 112.6 48.96 via_1600x480 ;
      VIA 92.4 48.96 via3_1600x480 ;
      VIA 92.4 48.96 via2_1600x480 ;
      VIA 92.4 48.96 via_1600x480 ;
      VIA 72.2 48.96 via3_1600x480 ;
      VIA 72.2 48.96 via2_1600x480 ;
      VIA 72.2 48.96 via_1600x480 ;
      VIA 52 48.96 via3_1600x480 ;
      VIA 52 48.96 via2_1600x480 ;
      VIA 52 48.96 via_1600x480 ;
      VIA 31.8 48.96 via3_1600x480 ;
      VIA 31.8 48.96 via2_1600x480 ;
      VIA 31.8 48.96 via_1600x480 ;
      VIA 11.6 48.96 via3_1600x480 ;
      VIA 11.6 48.96 via2_1600x480 ;
      VIA 11.6 48.96 via_1600x480 ;
      VIA 334.8 43.52 via3_1600x480 ;
      VIA 334.8 43.52 via2_1600x480 ;
      VIA 334.8 43.52 via_1600x480 ;
      VIA 314.6 43.52 via3_1600x480 ;
      VIA 314.6 43.52 via2_1600x480 ;
      VIA 314.6 43.52 via_1600x480 ;
      VIA 294.4 43.52 via3_1600x480 ;
      VIA 294.4 43.52 via2_1600x480 ;
      VIA 294.4 43.52 via_1600x480 ;
      VIA 274.2 43.52 via3_1600x480 ;
      VIA 274.2 43.52 via2_1600x480 ;
      VIA 274.2 43.52 via_1600x480 ;
      VIA 254 43.52 via3_1600x480 ;
      VIA 254 43.52 via2_1600x480 ;
      VIA 254 43.52 via_1600x480 ;
      VIA 233.8 43.52 via3_1600x480 ;
      VIA 233.8 43.52 via2_1600x480 ;
      VIA 233.8 43.52 via_1600x480 ;
      VIA 213.6 43.52 via3_1600x480 ;
      VIA 213.6 43.52 via2_1600x480 ;
      VIA 213.6 43.52 via_1600x480 ;
      VIA 193.4 43.52 via3_1600x480 ;
      VIA 193.4 43.52 via2_1600x480 ;
      VIA 193.4 43.52 via_1600x480 ;
      VIA 173.2 43.52 via3_1600x480 ;
      VIA 173.2 43.52 via2_1600x480 ;
      VIA 173.2 43.52 via_1600x480 ;
      VIA 153 43.52 via3_1600x480 ;
      VIA 153 43.52 via2_1600x480 ;
      VIA 153 43.52 via_1600x480 ;
      VIA 132.8 43.52 via3_1600x480 ;
      VIA 132.8 43.52 via2_1600x480 ;
      VIA 132.8 43.52 via_1600x480 ;
      VIA 112.6 43.52 via3_1600x480 ;
      VIA 112.6 43.52 via2_1600x480 ;
      VIA 112.6 43.52 via_1600x480 ;
      VIA 92.4 43.52 via3_1600x480 ;
      VIA 92.4 43.52 via2_1600x480 ;
      VIA 92.4 43.52 via_1600x480 ;
      VIA 72.2 43.52 via3_1600x480 ;
      VIA 72.2 43.52 via2_1600x480 ;
      VIA 72.2 43.52 via_1600x480 ;
      VIA 52 43.52 via3_1600x480 ;
      VIA 52 43.52 via2_1600x480 ;
      VIA 52 43.52 via_1600x480 ;
      VIA 31.8 43.52 via3_1600x480 ;
      VIA 31.8 43.52 via2_1600x480 ;
      VIA 31.8 43.52 via_1600x480 ;
      VIA 11.6 43.52 via3_1600x480 ;
      VIA 11.6 43.52 via2_1600x480 ;
      VIA 11.6 43.52 via_1600x480 ;
      VIA 334.8 38.08 via3_1600x480 ;
      VIA 334.8 38.08 via2_1600x480 ;
      VIA 334.8 38.08 via_1600x480 ;
      VIA 314.6 38.08 via3_1600x480 ;
      VIA 314.6 38.08 via2_1600x480 ;
      VIA 314.6 38.08 via_1600x480 ;
      VIA 294.4 38.08 via3_1600x480 ;
      VIA 294.4 38.08 via2_1600x480 ;
      VIA 294.4 38.08 via_1600x480 ;
      VIA 274.2 38.08 via3_1600x480 ;
      VIA 274.2 38.08 via2_1600x480 ;
      VIA 274.2 38.08 via_1600x480 ;
      VIA 254 38.08 via3_1600x480 ;
      VIA 254 38.08 via2_1600x480 ;
      VIA 254 38.08 via_1600x480 ;
      VIA 233.8 38.08 via3_1600x480 ;
      VIA 233.8 38.08 via2_1600x480 ;
      VIA 233.8 38.08 via_1600x480 ;
      VIA 213.6 38.08 via3_1600x480 ;
      VIA 213.6 38.08 via2_1600x480 ;
      VIA 213.6 38.08 via_1600x480 ;
      VIA 193.4 38.08 via3_1600x480 ;
      VIA 193.4 38.08 via2_1600x480 ;
      VIA 193.4 38.08 via_1600x480 ;
      VIA 173.2 38.08 via3_1600x480 ;
      VIA 173.2 38.08 via2_1600x480 ;
      VIA 173.2 38.08 via_1600x480 ;
      VIA 153 38.08 via3_1600x480 ;
      VIA 153 38.08 via2_1600x480 ;
      VIA 153 38.08 via_1600x480 ;
      VIA 132.8 38.08 via3_1600x480 ;
      VIA 132.8 38.08 via2_1600x480 ;
      VIA 132.8 38.08 via_1600x480 ;
      VIA 112.6 38.08 via3_1600x480 ;
      VIA 112.6 38.08 via2_1600x480 ;
      VIA 112.6 38.08 via_1600x480 ;
      VIA 92.4 38.08 via3_1600x480 ;
      VIA 92.4 38.08 via2_1600x480 ;
      VIA 92.4 38.08 via_1600x480 ;
      VIA 72.2 38.08 via3_1600x480 ;
      VIA 72.2 38.08 via2_1600x480 ;
      VIA 72.2 38.08 via_1600x480 ;
      VIA 52 38.08 via3_1600x480 ;
      VIA 52 38.08 via2_1600x480 ;
      VIA 52 38.08 via_1600x480 ;
      VIA 31.8 38.08 via3_1600x480 ;
      VIA 31.8 38.08 via2_1600x480 ;
      VIA 31.8 38.08 via_1600x480 ;
      VIA 11.6 38.08 via3_1600x480 ;
      VIA 11.6 38.08 via2_1600x480 ;
      VIA 11.6 38.08 via_1600x480 ;
      VIA 334.8 32.64 via3_1600x480 ;
      VIA 334.8 32.64 via2_1600x480 ;
      VIA 334.8 32.64 via_1600x480 ;
      VIA 314.6 32.64 via3_1600x480 ;
      VIA 314.6 32.64 via2_1600x480 ;
      VIA 314.6 32.64 via_1600x480 ;
      VIA 294.4 32.64 via3_1600x480 ;
      VIA 294.4 32.64 via2_1600x480 ;
      VIA 294.4 32.64 via_1600x480 ;
      VIA 274.2 32.64 via3_1600x480 ;
      VIA 274.2 32.64 via2_1600x480 ;
      VIA 274.2 32.64 via_1600x480 ;
      VIA 254 32.64 via3_1600x480 ;
      VIA 254 32.64 via2_1600x480 ;
      VIA 254 32.64 via_1600x480 ;
      VIA 233.8 32.64 via3_1600x480 ;
      VIA 233.8 32.64 via2_1600x480 ;
      VIA 233.8 32.64 via_1600x480 ;
      VIA 213.6 32.64 via3_1600x480 ;
      VIA 213.6 32.64 via2_1600x480 ;
      VIA 213.6 32.64 via_1600x480 ;
      VIA 193.4 32.64 via3_1600x480 ;
      VIA 193.4 32.64 via2_1600x480 ;
      VIA 193.4 32.64 via_1600x480 ;
      VIA 173.2 32.64 via3_1600x480 ;
      VIA 173.2 32.64 via2_1600x480 ;
      VIA 173.2 32.64 via_1600x480 ;
      VIA 153 32.64 via3_1600x480 ;
      VIA 153 32.64 via2_1600x480 ;
      VIA 153 32.64 via_1600x480 ;
      VIA 132.8 32.64 via3_1600x480 ;
      VIA 132.8 32.64 via2_1600x480 ;
      VIA 132.8 32.64 via_1600x480 ;
      VIA 112.6 32.64 via3_1600x480 ;
      VIA 112.6 32.64 via2_1600x480 ;
      VIA 112.6 32.64 via_1600x480 ;
      VIA 92.4 32.64 via3_1600x480 ;
      VIA 92.4 32.64 via2_1600x480 ;
      VIA 92.4 32.64 via_1600x480 ;
      VIA 72.2 32.64 via3_1600x480 ;
      VIA 72.2 32.64 via2_1600x480 ;
      VIA 72.2 32.64 via_1600x480 ;
      VIA 52 32.64 via3_1600x480 ;
      VIA 52 32.64 via2_1600x480 ;
      VIA 52 32.64 via_1600x480 ;
      VIA 31.8 32.64 via3_1600x480 ;
      VIA 31.8 32.64 via2_1600x480 ;
      VIA 31.8 32.64 via_1600x480 ;
      VIA 11.6 32.64 via3_1600x480 ;
      VIA 11.6 32.64 via2_1600x480 ;
      VIA 11.6 32.64 via_1600x480 ;
      VIA 334.8 27.2 via3_1600x480 ;
      VIA 334.8 27.2 via2_1600x480 ;
      VIA 334.8 27.2 via_1600x480 ;
      VIA 314.6 27.2 via3_1600x480 ;
      VIA 314.6 27.2 via2_1600x480 ;
      VIA 314.6 27.2 via_1600x480 ;
      VIA 294.4 27.2 via3_1600x480 ;
      VIA 294.4 27.2 via2_1600x480 ;
      VIA 294.4 27.2 via_1600x480 ;
      VIA 274.2 27.2 via3_1600x480 ;
      VIA 274.2 27.2 via2_1600x480 ;
      VIA 274.2 27.2 via_1600x480 ;
      VIA 254 27.2 via3_1600x480 ;
      VIA 254 27.2 via2_1600x480 ;
      VIA 254 27.2 via_1600x480 ;
      VIA 233.8 27.2 via3_1600x480 ;
      VIA 233.8 27.2 via2_1600x480 ;
      VIA 233.8 27.2 via_1600x480 ;
      VIA 213.6 27.2 via3_1600x480 ;
      VIA 213.6 27.2 via2_1600x480 ;
      VIA 213.6 27.2 via_1600x480 ;
      VIA 193.4 27.2 via3_1600x480 ;
      VIA 193.4 27.2 via2_1600x480 ;
      VIA 193.4 27.2 via_1600x480 ;
      VIA 173.2 27.2 via3_1600x480 ;
      VIA 173.2 27.2 via2_1600x480 ;
      VIA 173.2 27.2 via_1600x480 ;
      VIA 153 27.2 via3_1600x480 ;
      VIA 153 27.2 via2_1600x480 ;
      VIA 153 27.2 via_1600x480 ;
      VIA 132.8 27.2 via3_1600x480 ;
      VIA 132.8 27.2 via2_1600x480 ;
      VIA 132.8 27.2 via_1600x480 ;
      VIA 112.6 27.2 via3_1600x480 ;
      VIA 112.6 27.2 via2_1600x480 ;
      VIA 112.6 27.2 via_1600x480 ;
      VIA 92.4 27.2 via3_1600x480 ;
      VIA 92.4 27.2 via2_1600x480 ;
      VIA 92.4 27.2 via_1600x480 ;
      VIA 72.2 27.2 via3_1600x480 ;
      VIA 72.2 27.2 via2_1600x480 ;
      VIA 72.2 27.2 via_1600x480 ;
      VIA 52 27.2 via3_1600x480 ;
      VIA 52 27.2 via2_1600x480 ;
      VIA 52 27.2 via_1600x480 ;
      VIA 31.8 27.2 via3_1600x480 ;
      VIA 31.8 27.2 via2_1600x480 ;
      VIA 31.8 27.2 via_1600x480 ;
      VIA 11.6 27.2 via3_1600x480 ;
      VIA 11.6 27.2 via2_1600x480 ;
      VIA 11.6 27.2 via_1600x480 ;
      VIA 334.8 21.76 via3_1600x480 ;
      VIA 334.8 21.76 via2_1600x480 ;
      VIA 334.8 21.76 via_1600x480 ;
      VIA 314.6 21.76 via3_1600x480 ;
      VIA 314.6 21.76 via2_1600x480 ;
      VIA 314.6 21.76 via_1600x480 ;
      VIA 294.4 21.76 via3_1600x480 ;
      VIA 294.4 21.76 via2_1600x480 ;
      VIA 294.4 21.76 via_1600x480 ;
      VIA 274.2 21.76 via3_1600x480 ;
      VIA 274.2 21.76 via2_1600x480 ;
      VIA 274.2 21.76 via_1600x480 ;
      VIA 254 21.76 via3_1600x480 ;
      VIA 254 21.76 via2_1600x480 ;
      VIA 254 21.76 via_1600x480 ;
      VIA 233.8 21.76 via3_1600x480 ;
      VIA 233.8 21.76 via2_1600x480 ;
      VIA 233.8 21.76 via_1600x480 ;
      VIA 213.6 21.76 via3_1600x480 ;
      VIA 213.6 21.76 via2_1600x480 ;
      VIA 213.6 21.76 via_1600x480 ;
      VIA 193.4 21.76 via3_1600x480 ;
      VIA 193.4 21.76 via2_1600x480 ;
      VIA 193.4 21.76 via_1600x480 ;
      VIA 173.2 21.76 via3_1600x480 ;
      VIA 173.2 21.76 via2_1600x480 ;
      VIA 173.2 21.76 via_1600x480 ;
      VIA 153 21.76 via3_1600x480 ;
      VIA 153 21.76 via2_1600x480 ;
      VIA 153 21.76 via_1600x480 ;
      VIA 132.8 21.76 via3_1600x480 ;
      VIA 132.8 21.76 via2_1600x480 ;
      VIA 132.8 21.76 via_1600x480 ;
      VIA 112.6 21.76 via3_1600x480 ;
      VIA 112.6 21.76 via2_1600x480 ;
      VIA 112.6 21.76 via_1600x480 ;
      VIA 92.4 21.76 via3_1600x480 ;
      VIA 92.4 21.76 via2_1600x480 ;
      VIA 92.4 21.76 via_1600x480 ;
      VIA 72.2 21.76 via3_1600x480 ;
      VIA 72.2 21.76 via2_1600x480 ;
      VIA 72.2 21.76 via_1600x480 ;
      VIA 52 21.76 via3_1600x480 ;
      VIA 52 21.76 via2_1600x480 ;
      VIA 52 21.76 via_1600x480 ;
      VIA 31.8 21.76 via3_1600x480 ;
      VIA 31.8 21.76 via2_1600x480 ;
      VIA 31.8 21.76 via_1600x480 ;
      VIA 11.6 21.76 via3_1600x480 ;
      VIA 11.6 21.76 via2_1600x480 ;
      VIA 11.6 21.76 via_1600x480 ;
      VIA 334.8 16.32 via3_1600x480 ;
      VIA 334.8 16.32 via2_1600x480 ;
      VIA 334.8 16.32 via_1600x480 ;
      VIA 314.6 16.32 via3_1600x480 ;
      VIA 314.6 16.32 via2_1600x480 ;
      VIA 314.6 16.32 via_1600x480 ;
      VIA 294.4 16.32 via3_1600x480 ;
      VIA 294.4 16.32 via2_1600x480 ;
      VIA 294.4 16.32 via_1600x480 ;
      VIA 274.2 16.32 via3_1600x480 ;
      VIA 274.2 16.32 via2_1600x480 ;
      VIA 274.2 16.32 via_1600x480 ;
      VIA 254 16.32 via3_1600x480 ;
      VIA 254 16.32 via2_1600x480 ;
      VIA 254 16.32 via_1600x480 ;
      VIA 233.8 16.32 via3_1600x480 ;
      VIA 233.8 16.32 via2_1600x480 ;
      VIA 233.8 16.32 via_1600x480 ;
      VIA 213.6 16.32 via3_1600x480 ;
      VIA 213.6 16.32 via2_1600x480 ;
      VIA 213.6 16.32 via_1600x480 ;
      VIA 193.4 16.32 via3_1600x480 ;
      VIA 193.4 16.32 via2_1600x480 ;
      VIA 193.4 16.32 via_1600x480 ;
      VIA 173.2 16.32 via3_1600x480 ;
      VIA 173.2 16.32 via2_1600x480 ;
      VIA 173.2 16.32 via_1600x480 ;
      VIA 153 16.32 via3_1600x480 ;
      VIA 153 16.32 via2_1600x480 ;
      VIA 153 16.32 via_1600x480 ;
      VIA 132.8 16.32 via3_1600x480 ;
      VIA 132.8 16.32 via2_1600x480 ;
      VIA 132.8 16.32 via_1600x480 ;
      VIA 112.6 16.32 via3_1600x480 ;
      VIA 112.6 16.32 via2_1600x480 ;
      VIA 112.6 16.32 via_1600x480 ;
      VIA 92.4 16.32 via3_1600x480 ;
      VIA 92.4 16.32 via2_1600x480 ;
      VIA 92.4 16.32 via_1600x480 ;
      VIA 72.2 16.32 via3_1600x480 ;
      VIA 72.2 16.32 via2_1600x480 ;
      VIA 72.2 16.32 via_1600x480 ;
      VIA 52 16.32 via3_1600x480 ;
      VIA 52 16.32 via2_1600x480 ;
      VIA 52 16.32 via_1600x480 ;
      VIA 31.8 16.32 via3_1600x480 ;
      VIA 31.8 16.32 via2_1600x480 ;
      VIA 31.8 16.32 via_1600x480 ;
      VIA 11.6 16.32 via3_1600x480 ;
      VIA 11.6 16.32 via2_1600x480 ;
      VIA 11.6 16.32 via_1600x480 ;
      VIA 334.8 10.88 via3_1600x480 ;
      VIA 334.8 10.88 via2_1600x480 ;
      VIA 334.8 10.88 via_1600x480 ;
      VIA 314.6 10.88 via3_1600x480 ;
      VIA 314.6 10.88 via2_1600x480 ;
      VIA 314.6 10.88 via_1600x480 ;
      VIA 294.4 10.88 via3_1600x480 ;
      VIA 294.4 10.88 via2_1600x480 ;
      VIA 294.4 10.88 via_1600x480 ;
      VIA 274.2 10.88 via3_1600x480 ;
      VIA 274.2 10.88 via2_1600x480 ;
      VIA 274.2 10.88 via_1600x480 ;
      VIA 254 10.88 via3_1600x480 ;
      VIA 254 10.88 via2_1600x480 ;
      VIA 254 10.88 via_1600x480 ;
      VIA 233.8 10.88 via3_1600x480 ;
      VIA 233.8 10.88 via2_1600x480 ;
      VIA 233.8 10.88 via_1600x480 ;
      VIA 213.6 10.88 via3_1600x480 ;
      VIA 213.6 10.88 via2_1600x480 ;
      VIA 213.6 10.88 via_1600x480 ;
      VIA 193.4 10.88 via3_1600x480 ;
      VIA 193.4 10.88 via2_1600x480 ;
      VIA 193.4 10.88 via_1600x480 ;
      VIA 173.2 10.88 via3_1600x480 ;
      VIA 173.2 10.88 via2_1600x480 ;
      VIA 173.2 10.88 via_1600x480 ;
      VIA 153 10.88 via3_1600x480 ;
      VIA 153 10.88 via2_1600x480 ;
      VIA 153 10.88 via_1600x480 ;
      VIA 132.8 10.88 via3_1600x480 ;
      VIA 132.8 10.88 via2_1600x480 ;
      VIA 132.8 10.88 via_1600x480 ;
      VIA 112.6 10.88 via3_1600x480 ;
      VIA 112.6 10.88 via2_1600x480 ;
      VIA 112.6 10.88 via_1600x480 ;
      VIA 92.4 10.88 via3_1600x480 ;
      VIA 92.4 10.88 via2_1600x480 ;
      VIA 92.4 10.88 via_1600x480 ;
      VIA 72.2 10.88 via3_1600x480 ;
      VIA 72.2 10.88 via2_1600x480 ;
      VIA 72.2 10.88 via_1600x480 ;
      VIA 52 10.88 via3_1600x480 ;
      VIA 52 10.88 via2_1600x480 ;
      VIA 52 10.88 via_1600x480 ;
      VIA 31.8 10.88 via3_1600x480 ;
      VIA 31.8 10.88 via2_1600x480 ;
      VIA 31.8 10.88 via_1600x480 ;
      VIA 11.6 10.88 via3_1600x480 ;
      VIA 11.6 10.88 via2_1600x480 ;
      VIA 11.6 10.88 via_1600x480 ;
      VIA 334.8 5.44 via3_1600x480 ;
      VIA 334.8 5.44 via2_1600x480 ;
      VIA 334.8 5.44 via_1600x480 ;
      VIA 314.6 5.44 via3_1600x480 ;
      VIA 314.6 5.44 via2_1600x480 ;
      VIA 314.6 5.44 via_1600x480 ;
      VIA 294.4 5.44 via3_1600x480 ;
      VIA 294.4 5.44 via2_1600x480 ;
      VIA 294.4 5.44 via_1600x480 ;
      VIA 274.2 5.44 via3_1600x480 ;
      VIA 274.2 5.44 via2_1600x480 ;
      VIA 274.2 5.44 via_1600x480 ;
      VIA 254 5.44 via3_1600x480 ;
      VIA 254 5.44 via2_1600x480 ;
      VIA 254 5.44 via_1600x480 ;
      VIA 233.8 5.44 via3_1600x480 ;
      VIA 233.8 5.44 via2_1600x480 ;
      VIA 233.8 5.44 via_1600x480 ;
      VIA 213.6 5.44 via3_1600x480 ;
      VIA 213.6 5.44 via2_1600x480 ;
      VIA 213.6 5.44 via_1600x480 ;
      VIA 193.4 5.44 via3_1600x480 ;
      VIA 193.4 5.44 via2_1600x480 ;
      VIA 193.4 5.44 via_1600x480 ;
      VIA 173.2 5.44 via3_1600x480 ;
      VIA 173.2 5.44 via2_1600x480 ;
      VIA 173.2 5.44 via_1600x480 ;
      VIA 153 5.44 via3_1600x480 ;
      VIA 153 5.44 via2_1600x480 ;
      VIA 153 5.44 via_1600x480 ;
      VIA 132.8 5.44 via3_1600x480 ;
      VIA 132.8 5.44 via2_1600x480 ;
      VIA 132.8 5.44 via_1600x480 ;
      VIA 112.6 5.44 via3_1600x480 ;
      VIA 112.6 5.44 via2_1600x480 ;
      VIA 112.6 5.44 via_1600x480 ;
      VIA 92.4 5.44 via3_1600x480 ;
      VIA 92.4 5.44 via2_1600x480 ;
      VIA 92.4 5.44 via_1600x480 ;
      VIA 72.2 5.44 via3_1600x480 ;
      VIA 72.2 5.44 via2_1600x480 ;
      VIA 72.2 5.44 via_1600x480 ;
      VIA 52 5.44 via3_1600x480 ;
      VIA 52 5.44 via2_1600x480 ;
      VIA 52 5.44 via_1600x480 ;
      VIA 31.8 5.44 via3_1600x480 ;
      VIA 31.8 5.44 via2_1600x480 ;
      VIA 31.8 5.44 via_1600x480 ;
      VIA 11.6 5.44 via3_1600x480 ;
      VIA 11.6 5.44 via2_1600x480 ;
      VIA 11.6 5.44 via_1600x480 ;
      LAYER met5 ;
        RECT  0 195.08 349.6 196.68 ;
        RECT  0 174.88 349.6 176.48 ;
        RECT  0 154.68 349.6 156.28 ;
        RECT  0 134.48 349.6 136.08 ;
        RECT  0 114.28 349.6 115.88 ;
        RECT  0 94.08 349.6 95.68 ;
        RECT  0 73.88 349.6 75.48 ;
        RECT  0 53.68 349.6 55.28 ;
        RECT  0 33.48 349.6 35.08 ;
        RECT  0 13.28 349.6 14.88 ;
      LAYER met4 ;
        RECT  334 2.48 335.6 198.8 ;
        RECT  313.8 2.48 315.4 198.8 ;
        RECT  293.6 2.48 295.2 198.8 ;
        RECT  273.4 2.48 275 198.8 ;
        RECT  253.2 2.48 254.8 198.8 ;
        RECT  233 2.48 234.6 198.8 ;
        RECT  212.8 2.48 214.4 198.8 ;
        RECT  192.6 2.48 194.2 198.8 ;
        RECT  172.4 2.48 174 198.8 ;
        RECT  152.2 2.48 153.8 198.8 ;
        RECT  132 2.48 133.6 198.8 ;
        RECT  111.8 2.48 113.4 198.8 ;
        RECT  91.6 2.48 93.2 198.8 ;
        RECT  71.4 2.48 73 198.8 ;
        RECT  51.2 2.48 52.8 198.8 ;
        RECT  31 2.48 32.6 198.8 ;
        RECT  10.8 2.48 12.4 198.8 ;
      LAYER met1 ;
        RECT  0 195.6 349.6 196.08 ;
        RECT  0 190.16 349.6 190.64 ;
        RECT  0 184.72 349.6 185.2 ;
        RECT  0 179.28 349.6 179.76 ;
        RECT  0 173.84 349.6 174.32 ;
        RECT  0 168.4 349.6 168.88 ;
        RECT  0 162.96 349.6 163.44 ;
        RECT  0 157.52 349.6 158 ;
        RECT  0 152.08 349.6 152.56 ;
        RECT  0 146.64 349.6 147.12 ;
        RECT  0 141.2 349.6 141.68 ;
        RECT  0 135.76 349.6 136.24 ;
        RECT  0 130.32 349.6 130.8 ;
        RECT  0 124.88 349.6 125.36 ;
        RECT  0 119.44 349.6 119.92 ;
        RECT  0 114 349.6 114.48 ;
        RECT  0 108.56 349.6 109.04 ;
        RECT  0 103.12 349.6 103.6 ;
        RECT  0 97.68 349.6 98.16 ;
        RECT  0 92.24 349.6 92.72 ;
        RECT  0 86.8 349.6 87.28 ;
        RECT  0 81.36 349.6 81.84 ;
        RECT  0 75.92 349.6 76.4 ;
        RECT  0 70.48 349.6 70.96 ;
        RECT  0 65.04 349.6 65.52 ;
        RECT  0 59.6 349.6 60.08 ;
        RECT  0 54.16 349.6 54.64 ;
        RECT  0 48.72 349.6 49.2 ;
        RECT  0 43.28 349.6 43.76 ;
        RECT  0 37.84 349.6 38.32 ;
        RECT  0 32.4 349.6 32.88 ;
        RECT  0 26.96 349.6 27.44 ;
        RECT  0 21.52 349.6 22 ;
        RECT  0 16.08 349.6 16.56 ;
        RECT  0 10.64 349.6 11.12 ;
        RECT  0 5.2 349.6 5.68 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      VIA 344.9 185.78 via4_1600x1600 ;
      VIA 324.7 185.78 via4_1600x1600 ;
      VIA 304.5 185.78 via4_1600x1600 ;
      VIA 284.3 185.78 via4_1600x1600 ;
      VIA 264.1 185.78 via4_1600x1600 ;
      VIA 243.9 185.78 via4_1600x1600 ;
      VIA 223.7 185.78 via4_1600x1600 ;
      VIA 203.5 185.78 via4_1600x1600 ;
      VIA 183.3 185.78 via4_1600x1600 ;
      VIA 163.1 185.78 via4_1600x1600 ;
      VIA 142.9 185.78 via4_1600x1600 ;
      VIA 122.7 185.78 via4_1600x1600 ;
      VIA 102.5 185.78 via4_1600x1600 ;
      VIA 82.3 185.78 via4_1600x1600 ;
      VIA 62.1 185.78 via4_1600x1600 ;
      VIA 41.9 185.78 via4_1600x1600 ;
      VIA 21.7 185.78 via4_1600x1600 ;
      VIA 344.9 165.58 via4_1600x1600 ;
      VIA 324.7 165.58 via4_1600x1600 ;
      VIA 304.5 165.58 via4_1600x1600 ;
      VIA 284.3 165.58 via4_1600x1600 ;
      VIA 264.1 165.58 via4_1600x1600 ;
      VIA 243.9 165.58 via4_1600x1600 ;
      VIA 223.7 165.58 via4_1600x1600 ;
      VIA 203.5 165.58 via4_1600x1600 ;
      VIA 183.3 165.58 via4_1600x1600 ;
      VIA 163.1 165.58 via4_1600x1600 ;
      VIA 142.9 165.58 via4_1600x1600 ;
      VIA 122.7 165.58 via4_1600x1600 ;
      VIA 102.5 165.58 via4_1600x1600 ;
      VIA 82.3 165.58 via4_1600x1600 ;
      VIA 62.1 165.58 via4_1600x1600 ;
      VIA 41.9 165.58 via4_1600x1600 ;
      VIA 21.7 165.58 via4_1600x1600 ;
      VIA 344.9 145.38 via4_1600x1600 ;
      VIA 324.7 145.38 via4_1600x1600 ;
      VIA 304.5 145.38 via4_1600x1600 ;
      VIA 284.3 145.38 via4_1600x1600 ;
      VIA 264.1 145.38 via4_1600x1600 ;
      VIA 243.9 145.38 via4_1600x1600 ;
      VIA 223.7 145.38 via4_1600x1600 ;
      VIA 203.5 145.38 via4_1600x1600 ;
      VIA 183.3 145.38 via4_1600x1600 ;
      VIA 163.1 145.38 via4_1600x1600 ;
      VIA 142.9 145.38 via4_1600x1600 ;
      VIA 122.7 145.38 via4_1600x1600 ;
      VIA 102.5 145.38 via4_1600x1600 ;
      VIA 82.3 145.38 via4_1600x1600 ;
      VIA 62.1 145.38 via4_1600x1600 ;
      VIA 41.9 145.38 via4_1600x1600 ;
      VIA 21.7 145.38 via4_1600x1600 ;
      VIA 344.9 125.18 via4_1600x1600 ;
      VIA 324.7 125.18 via4_1600x1600 ;
      VIA 304.5 125.18 via4_1600x1600 ;
      VIA 284.3 125.18 via4_1600x1600 ;
      VIA 264.1 125.18 via4_1600x1600 ;
      VIA 243.9 125.18 via4_1600x1600 ;
      VIA 223.7 125.18 via4_1600x1600 ;
      VIA 203.5 125.18 via4_1600x1600 ;
      VIA 183.3 125.18 via4_1600x1600 ;
      VIA 163.1 125.18 via4_1600x1600 ;
      VIA 142.9 125.18 via4_1600x1600 ;
      VIA 122.7 125.18 via4_1600x1600 ;
      VIA 102.5 125.18 via4_1600x1600 ;
      VIA 82.3 125.18 via4_1600x1600 ;
      VIA 62.1 125.18 via4_1600x1600 ;
      VIA 41.9 125.18 via4_1600x1600 ;
      VIA 21.7 125.18 via4_1600x1600 ;
      VIA 344.9 104.98 via4_1600x1600 ;
      VIA 324.7 104.98 via4_1600x1600 ;
      VIA 304.5 104.98 via4_1600x1600 ;
      VIA 284.3 104.98 via4_1600x1600 ;
      VIA 264.1 104.98 via4_1600x1600 ;
      VIA 243.9 104.98 via4_1600x1600 ;
      VIA 223.7 104.98 via4_1600x1600 ;
      VIA 203.5 104.98 via4_1600x1600 ;
      VIA 183.3 104.98 via4_1600x1600 ;
      VIA 163.1 104.98 via4_1600x1600 ;
      VIA 142.9 104.98 via4_1600x1600 ;
      VIA 122.7 104.98 via4_1600x1600 ;
      VIA 102.5 104.98 via4_1600x1600 ;
      VIA 82.3 104.98 via4_1600x1600 ;
      VIA 62.1 104.98 via4_1600x1600 ;
      VIA 41.9 104.98 via4_1600x1600 ;
      VIA 21.7 104.98 via4_1600x1600 ;
      VIA 344.9 84.78 via4_1600x1600 ;
      VIA 324.7 84.78 via4_1600x1600 ;
      VIA 304.5 84.78 via4_1600x1600 ;
      VIA 284.3 84.78 via4_1600x1600 ;
      VIA 264.1 84.78 via4_1600x1600 ;
      VIA 243.9 84.78 via4_1600x1600 ;
      VIA 223.7 84.78 via4_1600x1600 ;
      VIA 203.5 84.78 via4_1600x1600 ;
      VIA 183.3 84.78 via4_1600x1600 ;
      VIA 163.1 84.78 via4_1600x1600 ;
      VIA 142.9 84.78 via4_1600x1600 ;
      VIA 122.7 84.78 via4_1600x1600 ;
      VIA 102.5 84.78 via4_1600x1600 ;
      VIA 82.3 84.78 via4_1600x1600 ;
      VIA 62.1 84.78 via4_1600x1600 ;
      VIA 41.9 84.78 via4_1600x1600 ;
      VIA 21.7 84.78 via4_1600x1600 ;
      VIA 344.9 64.58 via4_1600x1600 ;
      VIA 324.7 64.58 via4_1600x1600 ;
      VIA 304.5 64.58 via4_1600x1600 ;
      VIA 284.3 64.58 via4_1600x1600 ;
      VIA 264.1 64.58 via4_1600x1600 ;
      VIA 243.9 64.58 via4_1600x1600 ;
      VIA 223.7 64.58 via4_1600x1600 ;
      VIA 203.5 64.58 via4_1600x1600 ;
      VIA 183.3 64.58 via4_1600x1600 ;
      VIA 163.1 64.58 via4_1600x1600 ;
      VIA 142.9 64.58 via4_1600x1600 ;
      VIA 122.7 64.58 via4_1600x1600 ;
      VIA 102.5 64.58 via4_1600x1600 ;
      VIA 82.3 64.58 via4_1600x1600 ;
      VIA 62.1 64.58 via4_1600x1600 ;
      VIA 41.9 64.58 via4_1600x1600 ;
      VIA 21.7 64.58 via4_1600x1600 ;
      VIA 344.9 44.38 via4_1600x1600 ;
      VIA 324.7 44.38 via4_1600x1600 ;
      VIA 304.5 44.38 via4_1600x1600 ;
      VIA 284.3 44.38 via4_1600x1600 ;
      VIA 264.1 44.38 via4_1600x1600 ;
      VIA 243.9 44.38 via4_1600x1600 ;
      VIA 223.7 44.38 via4_1600x1600 ;
      VIA 203.5 44.38 via4_1600x1600 ;
      VIA 183.3 44.38 via4_1600x1600 ;
      VIA 163.1 44.38 via4_1600x1600 ;
      VIA 142.9 44.38 via4_1600x1600 ;
      VIA 122.7 44.38 via4_1600x1600 ;
      VIA 102.5 44.38 via4_1600x1600 ;
      VIA 82.3 44.38 via4_1600x1600 ;
      VIA 62.1 44.38 via4_1600x1600 ;
      VIA 41.9 44.38 via4_1600x1600 ;
      VIA 21.7 44.38 via4_1600x1600 ;
      VIA 344.9 24.18 via4_1600x1600 ;
      VIA 324.7 24.18 via4_1600x1600 ;
      VIA 304.5 24.18 via4_1600x1600 ;
      VIA 284.3 24.18 via4_1600x1600 ;
      VIA 264.1 24.18 via4_1600x1600 ;
      VIA 243.9 24.18 via4_1600x1600 ;
      VIA 223.7 24.18 via4_1600x1600 ;
      VIA 203.5 24.18 via4_1600x1600 ;
      VIA 183.3 24.18 via4_1600x1600 ;
      VIA 163.1 24.18 via4_1600x1600 ;
      VIA 142.9 24.18 via4_1600x1600 ;
      VIA 122.7 24.18 via4_1600x1600 ;
      VIA 102.5 24.18 via4_1600x1600 ;
      VIA 82.3 24.18 via4_1600x1600 ;
      VIA 62.1 24.18 via4_1600x1600 ;
      VIA 41.9 24.18 via4_1600x1600 ;
      VIA 21.7 24.18 via4_1600x1600 ;
      VIA 344.9 198.56 via3_1600x480 ;
      VIA 344.9 198.56 via2_1600x480 ;
      VIA 344.9 198.56 via_1600x480 ;
      VIA 324.7 198.56 via3_1600x480 ;
      VIA 324.7 198.56 via2_1600x480 ;
      VIA 324.7 198.56 via_1600x480 ;
      VIA 304.5 198.56 via3_1600x480 ;
      VIA 304.5 198.56 via2_1600x480 ;
      VIA 304.5 198.56 via_1600x480 ;
      VIA 284.3 198.56 via3_1600x480 ;
      VIA 284.3 198.56 via2_1600x480 ;
      VIA 284.3 198.56 via_1600x480 ;
      VIA 264.1 198.56 via3_1600x480 ;
      VIA 264.1 198.56 via2_1600x480 ;
      VIA 264.1 198.56 via_1600x480 ;
      VIA 243.9 198.56 via3_1600x480 ;
      VIA 243.9 198.56 via2_1600x480 ;
      VIA 243.9 198.56 via_1600x480 ;
      VIA 223.7 198.56 via3_1600x480 ;
      VIA 223.7 198.56 via2_1600x480 ;
      VIA 223.7 198.56 via_1600x480 ;
      VIA 203.5 198.56 via3_1600x480 ;
      VIA 203.5 198.56 via2_1600x480 ;
      VIA 203.5 198.56 via_1600x480 ;
      VIA 183.3 198.56 via3_1600x480 ;
      VIA 183.3 198.56 via2_1600x480 ;
      VIA 183.3 198.56 via_1600x480 ;
      VIA 163.1 198.56 via3_1600x480 ;
      VIA 163.1 198.56 via2_1600x480 ;
      VIA 163.1 198.56 via_1600x480 ;
      VIA 142.9 198.56 via3_1600x480 ;
      VIA 142.9 198.56 via2_1600x480 ;
      VIA 142.9 198.56 via_1600x480 ;
      VIA 122.7 198.56 via3_1600x480 ;
      VIA 122.7 198.56 via2_1600x480 ;
      VIA 122.7 198.56 via_1600x480 ;
      VIA 102.5 198.56 via3_1600x480 ;
      VIA 102.5 198.56 via2_1600x480 ;
      VIA 102.5 198.56 via_1600x480 ;
      VIA 82.3 198.56 via3_1600x480 ;
      VIA 82.3 198.56 via2_1600x480 ;
      VIA 82.3 198.56 via_1600x480 ;
      VIA 62.1 198.56 via3_1600x480 ;
      VIA 62.1 198.56 via2_1600x480 ;
      VIA 62.1 198.56 via_1600x480 ;
      VIA 41.9 198.56 via3_1600x480 ;
      VIA 41.9 198.56 via2_1600x480 ;
      VIA 41.9 198.56 via_1600x480 ;
      VIA 21.7 198.56 via3_1600x480 ;
      VIA 21.7 198.56 via2_1600x480 ;
      VIA 21.7 198.56 via_1600x480 ;
      VIA 344.9 193.12 via3_1600x480 ;
      VIA 344.9 193.12 via2_1600x480 ;
      VIA 344.9 193.12 via_1600x480 ;
      VIA 324.7 193.12 via3_1600x480 ;
      VIA 324.7 193.12 via2_1600x480 ;
      VIA 324.7 193.12 via_1600x480 ;
      VIA 304.5 193.12 via3_1600x480 ;
      VIA 304.5 193.12 via2_1600x480 ;
      VIA 304.5 193.12 via_1600x480 ;
      VIA 284.3 193.12 via3_1600x480 ;
      VIA 284.3 193.12 via2_1600x480 ;
      VIA 284.3 193.12 via_1600x480 ;
      VIA 264.1 193.12 via3_1600x480 ;
      VIA 264.1 193.12 via2_1600x480 ;
      VIA 264.1 193.12 via_1600x480 ;
      VIA 243.9 193.12 via3_1600x480 ;
      VIA 243.9 193.12 via2_1600x480 ;
      VIA 243.9 193.12 via_1600x480 ;
      VIA 223.7 193.12 via3_1600x480 ;
      VIA 223.7 193.12 via2_1600x480 ;
      VIA 223.7 193.12 via_1600x480 ;
      VIA 203.5 193.12 via3_1600x480 ;
      VIA 203.5 193.12 via2_1600x480 ;
      VIA 203.5 193.12 via_1600x480 ;
      VIA 183.3 193.12 via3_1600x480 ;
      VIA 183.3 193.12 via2_1600x480 ;
      VIA 183.3 193.12 via_1600x480 ;
      VIA 163.1 193.12 via3_1600x480 ;
      VIA 163.1 193.12 via2_1600x480 ;
      VIA 163.1 193.12 via_1600x480 ;
      VIA 142.9 193.12 via3_1600x480 ;
      VIA 142.9 193.12 via2_1600x480 ;
      VIA 142.9 193.12 via_1600x480 ;
      VIA 122.7 193.12 via3_1600x480 ;
      VIA 122.7 193.12 via2_1600x480 ;
      VIA 122.7 193.12 via_1600x480 ;
      VIA 102.5 193.12 via3_1600x480 ;
      VIA 102.5 193.12 via2_1600x480 ;
      VIA 102.5 193.12 via_1600x480 ;
      VIA 82.3 193.12 via3_1600x480 ;
      VIA 82.3 193.12 via2_1600x480 ;
      VIA 82.3 193.12 via_1600x480 ;
      VIA 62.1 193.12 via3_1600x480 ;
      VIA 62.1 193.12 via2_1600x480 ;
      VIA 62.1 193.12 via_1600x480 ;
      VIA 41.9 193.12 via3_1600x480 ;
      VIA 41.9 193.12 via2_1600x480 ;
      VIA 41.9 193.12 via_1600x480 ;
      VIA 21.7 193.12 via3_1600x480 ;
      VIA 21.7 193.12 via2_1600x480 ;
      VIA 21.7 193.12 via_1600x480 ;
      VIA 344.9 187.68 via3_1600x480 ;
      VIA 344.9 187.68 via2_1600x480 ;
      VIA 344.9 187.68 via_1600x480 ;
      VIA 324.7 187.68 via3_1600x480 ;
      VIA 324.7 187.68 via2_1600x480 ;
      VIA 324.7 187.68 via_1600x480 ;
      VIA 304.5 187.68 via3_1600x480 ;
      VIA 304.5 187.68 via2_1600x480 ;
      VIA 304.5 187.68 via_1600x480 ;
      VIA 284.3 187.68 via3_1600x480 ;
      VIA 284.3 187.68 via2_1600x480 ;
      VIA 284.3 187.68 via_1600x480 ;
      VIA 264.1 187.68 via3_1600x480 ;
      VIA 264.1 187.68 via2_1600x480 ;
      VIA 264.1 187.68 via_1600x480 ;
      VIA 243.9 187.68 via3_1600x480 ;
      VIA 243.9 187.68 via2_1600x480 ;
      VIA 243.9 187.68 via_1600x480 ;
      VIA 223.7 187.68 via3_1600x480 ;
      VIA 223.7 187.68 via2_1600x480 ;
      VIA 223.7 187.68 via_1600x480 ;
      VIA 203.5 187.68 via3_1600x480 ;
      VIA 203.5 187.68 via2_1600x480 ;
      VIA 203.5 187.68 via_1600x480 ;
      VIA 183.3 187.68 via3_1600x480 ;
      VIA 183.3 187.68 via2_1600x480 ;
      VIA 183.3 187.68 via_1600x480 ;
      VIA 163.1 187.68 via3_1600x480 ;
      VIA 163.1 187.68 via2_1600x480 ;
      VIA 163.1 187.68 via_1600x480 ;
      VIA 142.9 187.68 via3_1600x480 ;
      VIA 142.9 187.68 via2_1600x480 ;
      VIA 142.9 187.68 via_1600x480 ;
      VIA 122.7 187.68 via3_1600x480 ;
      VIA 122.7 187.68 via2_1600x480 ;
      VIA 122.7 187.68 via_1600x480 ;
      VIA 102.5 187.68 via3_1600x480 ;
      VIA 102.5 187.68 via2_1600x480 ;
      VIA 102.5 187.68 via_1600x480 ;
      VIA 82.3 187.68 via3_1600x480 ;
      VIA 82.3 187.68 via2_1600x480 ;
      VIA 82.3 187.68 via_1600x480 ;
      VIA 62.1 187.68 via3_1600x480 ;
      VIA 62.1 187.68 via2_1600x480 ;
      VIA 62.1 187.68 via_1600x480 ;
      VIA 41.9 187.68 via3_1600x480 ;
      VIA 41.9 187.68 via2_1600x480 ;
      VIA 41.9 187.68 via_1600x480 ;
      VIA 21.7 187.68 via3_1600x480 ;
      VIA 21.7 187.68 via2_1600x480 ;
      VIA 21.7 187.68 via_1600x480 ;
      VIA 344.9 182.24 via3_1600x480 ;
      VIA 344.9 182.24 via2_1600x480 ;
      VIA 344.9 182.24 via_1600x480 ;
      VIA 324.7 182.24 via3_1600x480 ;
      VIA 324.7 182.24 via2_1600x480 ;
      VIA 324.7 182.24 via_1600x480 ;
      VIA 304.5 182.24 via3_1600x480 ;
      VIA 304.5 182.24 via2_1600x480 ;
      VIA 304.5 182.24 via_1600x480 ;
      VIA 284.3 182.24 via3_1600x480 ;
      VIA 284.3 182.24 via2_1600x480 ;
      VIA 284.3 182.24 via_1600x480 ;
      VIA 264.1 182.24 via3_1600x480 ;
      VIA 264.1 182.24 via2_1600x480 ;
      VIA 264.1 182.24 via_1600x480 ;
      VIA 243.9 182.24 via3_1600x480 ;
      VIA 243.9 182.24 via2_1600x480 ;
      VIA 243.9 182.24 via_1600x480 ;
      VIA 223.7 182.24 via3_1600x480 ;
      VIA 223.7 182.24 via2_1600x480 ;
      VIA 223.7 182.24 via_1600x480 ;
      VIA 203.5 182.24 via3_1600x480 ;
      VIA 203.5 182.24 via2_1600x480 ;
      VIA 203.5 182.24 via_1600x480 ;
      VIA 183.3 182.24 via3_1600x480 ;
      VIA 183.3 182.24 via2_1600x480 ;
      VIA 183.3 182.24 via_1600x480 ;
      VIA 163.1 182.24 via3_1600x480 ;
      VIA 163.1 182.24 via2_1600x480 ;
      VIA 163.1 182.24 via_1600x480 ;
      VIA 142.9 182.24 via3_1600x480 ;
      VIA 142.9 182.24 via2_1600x480 ;
      VIA 142.9 182.24 via_1600x480 ;
      VIA 122.7 182.24 via3_1600x480 ;
      VIA 122.7 182.24 via2_1600x480 ;
      VIA 122.7 182.24 via_1600x480 ;
      VIA 102.5 182.24 via3_1600x480 ;
      VIA 102.5 182.24 via2_1600x480 ;
      VIA 102.5 182.24 via_1600x480 ;
      VIA 82.3 182.24 via3_1600x480 ;
      VIA 82.3 182.24 via2_1600x480 ;
      VIA 82.3 182.24 via_1600x480 ;
      VIA 62.1 182.24 via3_1600x480 ;
      VIA 62.1 182.24 via2_1600x480 ;
      VIA 62.1 182.24 via_1600x480 ;
      VIA 41.9 182.24 via3_1600x480 ;
      VIA 41.9 182.24 via2_1600x480 ;
      VIA 41.9 182.24 via_1600x480 ;
      VIA 21.7 182.24 via3_1600x480 ;
      VIA 21.7 182.24 via2_1600x480 ;
      VIA 21.7 182.24 via_1600x480 ;
      VIA 344.9 176.8 via3_1600x480 ;
      VIA 344.9 176.8 via2_1600x480 ;
      VIA 344.9 176.8 via_1600x480 ;
      VIA 324.7 176.8 via3_1600x480 ;
      VIA 324.7 176.8 via2_1600x480 ;
      VIA 324.7 176.8 via_1600x480 ;
      VIA 304.5 176.8 via3_1600x480 ;
      VIA 304.5 176.8 via2_1600x480 ;
      VIA 304.5 176.8 via_1600x480 ;
      VIA 284.3 176.8 via3_1600x480 ;
      VIA 284.3 176.8 via2_1600x480 ;
      VIA 284.3 176.8 via_1600x480 ;
      VIA 264.1 176.8 via3_1600x480 ;
      VIA 264.1 176.8 via2_1600x480 ;
      VIA 264.1 176.8 via_1600x480 ;
      VIA 243.9 176.8 via3_1600x480 ;
      VIA 243.9 176.8 via2_1600x480 ;
      VIA 243.9 176.8 via_1600x480 ;
      VIA 223.7 176.8 via3_1600x480 ;
      VIA 223.7 176.8 via2_1600x480 ;
      VIA 223.7 176.8 via_1600x480 ;
      VIA 203.5 176.8 via3_1600x480 ;
      VIA 203.5 176.8 via2_1600x480 ;
      VIA 203.5 176.8 via_1600x480 ;
      VIA 183.3 176.8 via3_1600x480 ;
      VIA 183.3 176.8 via2_1600x480 ;
      VIA 183.3 176.8 via_1600x480 ;
      VIA 163.1 176.8 via3_1600x480 ;
      VIA 163.1 176.8 via2_1600x480 ;
      VIA 163.1 176.8 via_1600x480 ;
      VIA 142.9 176.8 via3_1600x480 ;
      VIA 142.9 176.8 via2_1600x480 ;
      VIA 142.9 176.8 via_1600x480 ;
      VIA 122.7 176.8 via3_1600x480 ;
      VIA 122.7 176.8 via2_1600x480 ;
      VIA 122.7 176.8 via_1600x480 ;
      VIA 102.5 176.8 via3_1600x480 ;
      VIA 102.5 176.8 via2_1600x480 ;
      VIA 102.5 176.8 via_1600x480 ;
      VIA 82.3 176.8 via3_1600x480 ;
      VIA 82.3 176.8 via2_1600x480 ;
      VIA 82.3 176.8 via_1600x480 ;
      VIA 62.1 176.8 via3_1600x480 ;
      VIA 62.1 176.8 via2_1600x480 ;
      VIA 62.1 176.8 via_1600x480 ;
      VIA 41.9 176.8 via3_1600x480 ;
      VIA 41.9 176.8 via2_1600x480 ;
      VIA 41.9 176.8 via_1600x480 ;
      VIA 21.7 176.8 via3_1600x480 ;
      VIA 21.7 176.8 via2_1600x480 ;
      VIA 21.7 176.8 via_1600x480 ;
      VIA 344.9 171.36 via3_1600x480 ;
      VIA 344.9 171.36 via2_1600x480 ;
      VIA 344.9 171.36 via_1600x480 ;
      VIA 324.7 171.36 via3_1600x480 ;
      VIA 324.7 171.36 via2_1600x480 ;
      VIA 324.7 171.36 via_1600x480 ;
      VIA 304.5 171.36 via3_1600x480 ;
      VIA 304.5 171.36 via2_1600x480 ;
      VIA 304.5 171.36 via_1600x480 ;
      VIA 284.3 171.36 via3_1600x480 ;
      VIA 284.3 171.36 via2_1600x480 ;
      VIA 284.3 171.36 via_1600x480 ;
      VIA 264.1 171.36 via3_1600x480 ;
      VIA 264.1 171.36 via2_1600x480 ;
      VIA 264.1 171.36 via_1600x480 ;
      VIA 243.9 171.36 via3_1600x480 ;
      VIA 243.9 171.36 via2_1600x480 ;
      VIA 243.9 171.36 via_1600x480 ;
      VIA 223.7 171.36 via3_1600x480 ;
      VIA 223.7 171.36 via2_1600x480 ;
      VIA 223.7 171.36 via_1600x480 ;
      VIA 203.5 171.36 via3_1600x480 ;
      VIA 203.5 171.36 via2_1600x480 ;
      VIA 203.5 171.36 via_1600x480 ;
      VIA 183.3 171.36 via3_1600x480 ;
      VIA 183.3 171.36 via2_1600x480 ;
      VIA 183.3 171.36 via_1600x480 ;
      VIA 163.1 171.36 via3_1600x480 ;
      VIA 163.1 171.36 via2_1600x480 ;
      VIA 163.1 171.36 via_1600x480 ;
      VIA 142.9 171.36 via3_1600x480 ;
      VIA 142.9 171.36 via2_1600x480 ;
      VIA 142.9 171.36 via_1600x480 ;
      VIA 122.7 171.36 via3_1600x480 ;
      VIA 122.7 171.36 via2_1600x480 ;
      VIA 122.7 171.36 via_1600x480 ;
      VIA 102.5 171.36 via3_1600x480 ;
      VIA 102.5 171.36 via2_1600x480 ;
      VIA 102.5 171.36 via_1600x480 ;
      VIA 82.3 171.36 via3_1600x480 ;
      VIA 82.3 171.36 via2_1600x480 ;
      VIA 82.3 171.36 via_1600x480 ;
      VIA 62.1 171.36 via3_1600x480 ;
      VIA 62.1 171.36 via2_1600x480 ;
      VIA 62.1 171.36 via_1600x480 ;
      VIA 41.9 171.36 via3_1600x480 ;
      VIA 41.9 171.36 via2_1600x480 ;
      VIA 41.9 171.36 via_1600x480 ;
      VIA 21.7 171.36 via3_1600x480 ;
      VIA 21.7 171.36 via2_1600x480 ;
      VIA 21.7 171.36 via_1600x480 ;
      VIA 344.9 165.92 via3_1600x480 ;
      VIA 344.9 165.92 via2_1600x480 ;
      VIA 344.9 165.92 via_1600x480 ;
      VIA 324.7 165.92 via3_1600x480 ;
      VIA 324.7 165.92 via2_1600x480 ;
      VIA 324.7 165.92 via_1600x480 ;
      VIA 304.5 165.92 via3_1600x480 ;
      VIA 304.5 165.92 via2_1600x480 ;
      VIA 304.5 165.92 via_1600x480 ;
      VIA 284.3 165.92 via3_1600x480 ;
      VIA 284.3 165.92 via2_1600x480 ;
      VIA 284.3 165.92 via_1600x480 ;
      VIA 264.1 165.92 via3_1600x480 ;
      VIA 264.1 165.92 via2_1600x480 ;
      VIA 264.1 165.92 via_1600x480 ;
      VIA 243.9 165.92 via3_1600x480 ;
      VIA 243.9 165.92 via2_1600x480 ;
      VIA 243.9 165.92 via_1600x480 ;
      VIA 223.7 165.92 via3_1600x480 ;
      VIA 223.7 165.92 via2_1600x480 ;
      VIA 223.7 165.92 via_1600x480 ;
      VIA 203.5 165.92 via3_1600x480 ;
      VIA 203.5 165.92 via2_1600x480 ;
      VIA 203.5 165.92 via_1600x480 ;
      VIA 183.3 165.92 via3_1600x480 ;
      VIA 183.3 165.92 via2_1600x480 ;
      VIA 183.3 165.92 via_1600x480 ;
      VIA 163.1 165.92 via3_1600x480 ;
      VIA 163.1 165.92 via2_1600x480 ;
      VIA 163.1 165.92 via_1600x480 ;
      VIA 142.9 165.92 via3_1600x480 ;
      VIA 142.9 165.92 via2_1600x480 ;
      VIA 142.9 165.92 via_1600x480 ;
      VIA 122.7 165.92 via3_1600x480 ;
      VIA 122.7 165.92 via2_1600x480 ;
      VIA 122.7 165.92 via_1600x480 ;
      VIA 102.5 165.92 via3_1600x480 ;
      VIA 102.5 165.92 via2_1600x480 ;
      VIA 102.5 165.92 via_1600x480 ;
      VIA 82.3 165.92 via3_1600x480 ;
      VIA 82.3 165.92 via2_1600x480 ;
      VIA 82.3 165.92 via_1600x480 ;
      VIA 62.1 165.92 via3_1600x480 ;
      VIA 62.1 165.92 via2_1600x480 ;
      VIA 62.1 165.92 via_1600x480 ;
      VIA 41.9 165.92 via3_1600x480 ;
      VIA 41.9 165.92 via2_1600x480 ;
      VIA 41.9 165.92 via_1600x480 ;
      VIA 21.7 165.92 via3_1600x480 ;
      VIA 21.7 165.92 via2_1600x480 ;
      VIA 21.7 165.92 via_1600x480 ;
      VIA 344.9 160.48 via3_1600x480 ;
      VIA 344.9 160.48 via2_1600x480 ;
      VIA 344.9 160.48 via_1600x480 ;
      VIA 324.7 160.48 via3_1600x480 ;
      VIA 324.7 160.48 via2_1600x480 ;
      VIA 324.7 160.48 via_1600x480 ;
      VIA 304.5 160.48 via3_1600x480 ;
      VIA 304.5 160.48 via2_1600x480 ;
      VIA 304.5 160.48 via_1600x480 ;
      VIA 284.3 160.48 via3_1600x480 ;
      VIA 284.3 160.48 via2_1600x480 ;
      VIA 284.3 160.48 via_1600x480 ;
      VIA 264.1 160.48 via3_1600x480 ;
      VIA 264.1 160.48 via2_1600x480 ;
      VIA 264.1 160.48 via_1600x480 ;
      VIA 243.9 160.48 via3_1600x480 ;
      VIA 243.9 160.48 via2_1600x480 ;
      VIA 243.9 160.48 via_1600x480 ;
      VIA 223.7 160.48 via3_1600x480 ;
      VIA 223.7 160.48 via2_1600x480 ;
      VIA 223.7 160.48 via_1600x480 ;
      VIA 203.5 160.48 via3_1600x480 ;
      VIA 203.5 160.48 via2_1600x480 ;
      VIA 203.5 160.48 via_1600x480 ;
      VIA 183.3 160.48 via3_1600x480 ;
      VIA 183.3 160.48 via2_1600x480 ;
      VIA 183.3 160.48 via_1600x480 ;
      VIA 163.1 160.48 via3_1600x480 ;
      VIA 163.1 160.48 via2_1600x480 ;
      VIA 163.1 160.48 via_1600x480 ;
      VIA 142.9 160.48 via3_1600x480 ;
      VIA 142.9 160.48 via2_1600x480 ;
      VIA 142.9 160.48 via_1600x480 ;
      VIA 122.7 160.48 via3_1600x480 ;
      VIA 122.7 160.48 via2_1600x480 ;
      VIA 122.7 160.48 via_1600x480 ;
      VIA 102.5 160.48 via3_1600x480 ;
      VIA 102.5 160.48 via2_1600x480 ;
      VIA 102.5 160.48 via_1600x480 ;
      VIA 82.3 160.48 via3_1600x480 ;
      VIA 82.3 160.48 via2_1600x480 ;
      VIA 82.3 160.48 via_1600x480 ;
      VIA 62.1 160.48 via3_1600x480 ;
      VIA 62.1 160.48 via2_1600x480 ;
      VIA 62.1 160.48 via_1600x480 ;
      VIA 41.9 160.48 via3_1600x480 ;
      VIA 41.9 160.48 via2_1600x480 ;
      VIA 41.9 160.48 via_1600x480 ;
      VIA 21.7 160.48 via3_1600x480 ;
      VIA 21.7 160.48 via2_1600x480 ;
      VIA 21.7 160.48 via_1600x480 ;
      VIA 344.9 155.04 via3_1600x480 ;
      VIA 344.9 155.04 via2_1600x480 ;
      VIA 344.9 155.04 via_1600x480 ;
      VIA 324.7 155.04 via3_1600x480 ;
      VIA 324.7 155.04 via2_1600x480 ;
      VIA 324.7 155.04 via_1600x480 ;
      VIA 304.5 155.04 via3_1600x480 ;
      VIA 304.5 155.04 via2_1600x480 ;
      VIA 304.5 155.04 via_1600x480 ;
      VIA 284.3 155.04 via3_1600x480 ;
      VIA 284.3 155.04 via2_1600x480 ;
      VIA 284.3 155.04 via_1600x480 ;
      VIA 264.1 155.04 via3_1600x480 ;
      VIA 264.1 155.04 via2_1600x480 ;
      VIA 264.1 155.04 via_1600x480 ;
      VIA 243.9 155.04 via3_1600x480 ;
      VIA 243.9 155.04 via2_1600x480 ;
      VIA 243.9 155.04 via_1600x480 ;
      VIA 223.7 155.04 via3_1600x480 ;
      VIA 223.7 155.04 via2_1600x480 ;
      VIA 223.7 155.04 via_1600x480 ;
      VIA 203.5 155.04 via3_1600x480 ;
      VIA 203.5 155.04 via2_1600x480 ;
      VIA 203.5 155.04 via_1600x480 ;
      VIA 183.3 155.04 via3_1600x480 ;
      VIA 183.3 155.04 via2_1600x480 ;
      VIA 183.3 155.04 via_1600x480 ;
      VIA 163.1 155.04 via3_1600x480 ;
      VIA 163.1 155.04 via2_1600x480 ;
      VIA 163.1 155.04 via_1600x480 ;
      VIA 142.9 155.04 via3_1600x480 ;
      VIA 142.9 155.04 via2_1600x480 ;
      VIA 142.9 155.04 via_1600x480 ;
      VIA 122.7 155.04 via3_1600x480 ;
      VIA 122.7 155.04 via2_1600x480 ;
      VIA 122.7 155.04 via_1600x480 ;
      VIA 102.5 155.04 via3_1600x480 ;
      VIA 102.5 155.04 via2_1600x480 ;
      VIA 102.5 155.04 via_1600x480 ;
      VIA 82.3 155.04 via3_1600x480 ;
      VIA 82.3 155.04 via2_1600x480 ;
      VIA 82.3 155.04 via_1600x480 ;
      VIA 62.1 155.04 via3_1600x480 ;
      VIA 62.1 155.04 via2_1600x480 ;
      VIA 62.1 155.04 via_1600x480 ;
      VIA 41.9 155.04 via3_1600x480 ;
      VIA 41.9 155.04 via2_1600x480 ;
      VIA 41.9 155.04 via_1600x480 ;
      VIA 21.7 155.04 via3_1600x480 ;
      VIA 21.7 155.04 via2_1600x480 ;
      VIA 21.7 155.04 via_1600x480 ;
      VIA 344.9 149.6 via3_1600x480 ;
      VIA 344.9 149.6 via2_1600x480 ;
      VIA 344.9 149.6 via_1600x480 ;
      VIA 324.7 149.6 via3_1600x480 ;
      VIA 324.7 149.6 via2_1600x480 ;
      VIA 324.7 149.6 via_1600x480 ;
      VIA 304.5 149.6 via3_1600x480 ;
      VIA 304.5 149.6 via2_1600x480 ;
      VIA 304.5 149.6 via_1600x480 ;
      VIA 284.3 149.6 via3_1600x480 ;
      VIA 284.3 149.6 via2_1600x480 ;
      VIA 284.3 149.6 via_1600x480 ;
      VIA 264.1 149.6 via3_1600x480 ;
      VIA 264.1 149.6 via2_1600x480 ;
      VIA 264.1 149.6 via_1600x480 ;
      VIA 243.9 149.6 via3_1600x480 ;
      VIA 243.9 149.6 via2_1600x480 ;
      VIA 243.9 149.6 via_1600x480 ;
      VIA 223.7 149.6 via3_1600x480 ;
      VIA 223.7 149.6 via2_1600x480 ;
      VIA 223.7 149.6 via_1600x480 ;
      VIA 203.5 149.6 via3_1600x480 ;
      VIA 203.5 149.6 via2_1600x480 ;
      VIA 203.5 149.6 via_1600x480 ;
      VIA 183.3 149.6 via3_1600x480 ;
      VIA 183.3 149.6 via2_1600x480 ;
      VIA 183.3 149.6 via_1600x480 ;
      VIA 163.1 149.6 via3_1600x480 ;
      VIA 163.1 149.6 via2_1600x480 ;
      VIA 163.1 149.6 via_1600x480 ;
      VIA 142.9 149.6 via3_1600x480 ;
      VIA 142.9 149.6 via2_1600x480 ;
      VIA 142.9 149.6 via_1600x480 ;
      VIA 122.7 149.6 via3_1600x480 ;
      VIA 122.7 149.6 via2_1600x480 ;
      VIA 122.7 149.6 via_1600x480 ;
      VIA 102.5 149.6 via3_1600x480 ;
      VIA 102.5 149.6 via2_1600x480 ;
      VIA 102.5 149.6 via_1600x480 ;
      VIA 82.3 149.6 via3_1600x480 ;
      VIA 82.3 149.6 via2_1600x480 ;
      VIA 82.3 149.6 via_1600x480 ;
      VIA 62.1 149.6 via3_1600x480 ;
      VIA 62.1 149.6 via2_1600x480 ;
      VIA 62.1 149.6 via_1600x480 ;
      VIA 41.9 149.6 via3_1600x480 ;
      VIA 41.9 149.6 via2_1600x480 ;
      VIA 41.9 149.6 via_1600x480 ;
      VIA 21.7 149.6 via3_1600x480 ;
      VIA 21.7 149.6 via2_1600x480 ;
      VIA 21.7 149.6 via_1600x480 ;
      VIA 344.9 144.16 via3_1600x480 ;
      VIA 344.9 144.16 via2_1600x480 ;
      VIA 344.9 144.16 via_1600x480 ;
      VIA 324.7 144.16 via3_1600x480 ;
      VIA 324.7 144.16 via2_1600x480 ;
      VIA 324.7 144.16 via_1600x480 ;
      VIA 304.5 144.16 via3_1600x480 ;
      VIA 304.5 144.16 via2_1600x480 ;
      VIA 304.5 144.16 via_1600x480 ;
      VIA 284.3 144.16 via3_1600x480 ;
      VIA 284.3 144.16 via2_1600x480 ;
      VIA 284.3 144.16 via_1600x480 ;
      VIA 264.1 144.16 via3_1600x480 ;
      VIA 264.1 144.16 via2_1600x480 ;
      VIA 264.1 144.16 via_1600x480 ;
      VIA 243.9 144.16 via3_1600x480 ;
      VIA 243.9 144.16 via2_1600x480 ;
      VIA 243.9 144.16 via_1600x480 ;
      VIA 223.7 144.16 via3_1600x480 ;
      VIA 223.7 144.16 via2_1600x480 ;
      VIA 223.7 144.16 via_1600x480 ;
      VIA 203.5 144.16 via3_1600x480 ;
      VIA 203.5 144.16 via2_1600x480 ;
      VIA 203.5 144.16 via_1600x480 ;
      VIA 183.3 144.16 via3_1600x480 ;
      VIA 183.3 144.16 via2_1600x480 ;
      VIA 183.3 144.16 via_1600x480 ;
      VIA 163.1 144.16 via3_1600x480 ;
      VIA 163.1 144.16 via2_1600x480 ;
      VIA 163.1 144.16 via_1600x480 ;
      VIA 142.9 144.16 via3_1600x480 ;
      VIA 142.9 144.16 via2_1600x480 ;
      VIA 142.9 144.16 via_1600x480 ;
      VIA 122.7 144.16 via3_1600x480 ;
      VIA 122.7 144.16 via2_1600x480 ;
      VIA 122.7 144.16 via_1600x480 ;
      VIA 102.5 144.16 via3_1600x480 ;
      VIA 102.5 144.16 via2_1600x480 ;
      VIA 102.5 144.16 via_1600x480 ;
      VIA 82.3 144.16 via3_1600x480 ;
      VIA 82.3 144.16 via2_1600x480 ;
      VIA 82.3 144.16 via_1600x480 ;
      VIA 62.1 144.16 via3_1600x480 ;
      VIA 62.1 144.16 via2_1600x480 ;
      VIA 62.1 144.16 via_1600x480 ;
      VIA 41.9 144.16 via3_1600x480 ;
      VIA 41.9 144.16 via2_1600x480 ;
      VIA 41.9 144.16 via_1600x480 ;
      VIA 21.7 144.16 via3_1600x480 ;
      VIA 21.7 144.16 via2_1600x480 ;
      VIA 21.7 144.16 via_1600x480 ;
      VIA 344.9 138.72 via3_1600x480 ;
      VIA 344.9 138.72 via2_1600x480 ;
      VIA 344.9 138.72 via_1600x480 ;
      VIA 324.7 138.72 via3_1600x480 ;
      VIA 324.7 138.72 via2_1600x480 ;
      VIA 324.7 138.72 via_1600x480 ;
      VIA 304.5 138.72 via3_1600x480 ;
      VIA 304.5 138.72 via2_1600x480 ;
      VIA 304.5 138.72 via_1600x480 ;
      VIA 284.3 138.72 via3_1600x480 ;
      VIA 284.3 138.72 via2_1600x480 ;
      VIA 284.3 138.72 via_1600x480 ;
      VIA 264.1 138.72 via3_1600x480 ;
      VIA 264.1 138.72 via2_1600x480 ;
      VIA 264.1 138.72 via_1600x480 ;
      VIA 243.9 138.72 via3_1600x480 ;
      VIA 243.9 138.72 via2_1600x480 ;
      VIA 243.9 138.72 via_1600x480 ;
      VIA 223.7 138.72 via3_1600x480 ;
      VIA 223.7 138.72 via2_1600x480 ;
      VIA 223.7 138.72 via_1600x480 ;
      VIA 203.5 138.72 via3_1600x480 ;
      VIA 203.5 138.72 via2_1600x480 ;
      VIA 203.5 138.72 via_1600x480 ;
      VIA 183.3 138.72 via3_1600x480 ;
      VIA 183.3 138.72 via2_1600x480 ;
      VIA 183.3 138.72 via_1600x480 ;
      VIA 163.1 138.72 via3_1600x480 ;
      VIA 163.1 138.72 via2_1600x480 ;
      VIA 163.1 138.72 via_1600x480 ;
      VIA 142.9 138.72 via3_1600x480 ;
      VIA 142.9 138.72 via2_1600x480 ;
      VIA 142.9 138.72 via_1600x480 ;
      VIA 122.7 138.72 via3_1600x480 ;
      VIA 122.7 138.72 via2_1600x480 ;
      VIA 122.7 138.72 via_1600x480 ;
      VIA 102.5 138.72 via3_1600x480 ;
      VIA 102.5 138.72 via2_1600x480 ;
      VIA 102.5 138.72 via_1600x480 ;
      VIA 82.3 138.72 via3_1600x480 ;
      VIA 82.3 138.72 via2_1600x480 ;
      VIA 82.3 138.72 via_1600x480 ;
      VIA 62.1 138.72 via3_1600x480 ;
      VIA 62.1 138.72 via2_1600x480 ;
      VIA 62.1 138.72 via_1600x480 ;
      VIA 41.9 138.72 via3_1600x480 ;
      VIA 41.9 138.72 via2_1600x480 ;
      VIA 41.9 138.72 via_1600x480 ;
      VIA 21.7 138.72 via3_1600x480 ;
      VIA 21.7 138.72 via2_1600x480 ;
      VIA 21.7 138.72 via_1600x480 ;
      VIA 344.9 133.28 via3_1600x480 ;
      VIA 344.9 133.28 via2_1600x480 ;
      VIA 344.9 133.28 via_1600x480 ;
      VIA 324.7 133.28 via3_1600x480 ;
      VIA 324.7 133.28 via2_1600x480 ;
      VIA 324.7 133.28 via_1600x480 ;
      VIA 304.5 133.28 via3_1600x480 ;
      VIA 304.5 133.28 via2_1600x480 ;
      VIA 304.5 133.28 via_1600x480 ;
      VIA 284.3 133.28 via3_1600x480 ;
      VIA 284.3 133.28 via2_1600x480 ;
      VIA 284.3 133.28 via_1600x480 ;
      VIA 264.1 133.28 via3_1600x480 ;
      VIA 264.1 133.28 via2_1600x480 ;
      VIA 264.1 133.28 via_1600x480 ;
      VIA 243.9 133.28 via3_1600x480 ;
      VIA 243.9 133.28 via2_1600x480 ;
      VIA 243.9 133.28 via_1600x480 ;
      VIA 223.7 133.28 via3_1600x480 ;
      VIA 223.7 133.28 via2_1600x480 ;
      VIA 223.7 133.28 via_1600x480 ;
      VIA 203.5 133.28 via3_1600x480 ;
      VIA 203.5 133.28 via2_1600x480 ;
      VIA 203.5 133.28 via_1600x480 ;
      VIA 183.3 133.28 via3_1600x480 ;
      VIA 183.3 133.28 via2_1600x480 ;
      VIA 183.3 133.28 via_1600x480 ;
      VIA 163.1 133.28 via3_1600x480 ;
      VIA 163.1 133.28 via2_1600x480 ;
      VIA 163.1 133.28 via_1600x480 ;
      VIA 142.9 133.28 via3_1600x480 ;
      VIA 142.9 133.28 via2_1600x480 ;
      VIA 142.9 133.28 via_1600x480 ;
      VIA 122.7 133.28 via3_1600x480 ;
      VIA 122.7 133.28 via2_1600x480 ;
      VIA 122.7 133.28 via_1600x480 ;
      VIA 102.5 133.28 via3_1600x480 ;
      VIA 102.5 133.28 via2_1600x480 ;
      VIA 102.5 133.28 via_1600x480 ;
      VIA 82.3 133.28 via3_1600x480 ;
      VIA 82.3 133.28 via2_1600x480 ;
      VIA 82.3 133.28 via_1600x480 ;
      VIA 62.1 133.28 via3_1600x480 ;
      VIA 62.1 133.28 via2_1600x480 ;
      VIA 62.1 133.28 via_1600x480 ;
      VIA 41.9 133.28 via3_1600x480 ;
      VIA 41.9 133.28 via2_1600x480 ;
      VIA 41.9 133.28 via_1600x480 ;
      VIA 21.7 133.28 via3_1600x480 ;
      VIA 21.7 133.28 via2_1600x480 ;
      VIA 21.7 133.28 via_1600x480 ;
      VIA 344.9 127.84 via3_1600x480 ;
      VIA 344.9 127.84 via2_1600x480 ;
      VIA 344.9 127.84 via_1600x480 ;
      VIA 324.7 127.84 via3_1600x480 ;
      VIA 324.7 127.84 via2_1600x480 ;
      VIA 324.7 127.84 via_1600x480 ;
      VIA 304.5 127.84 via3_1600x480 ;
      VIA 304.5 127.84 via2_1600x480 ;
      VIA 304.5 127.84 via_1600x480 ;
      VIA 284.3 127.84 via3_1600x480 ;
      VIA 284.3 127.84 via2_1600x480 ;
      VIA 284.3 127.84 via_1600x480 ;
      VIA 264.1 127.84 via3_1600x480 ;
      VIA 264.1 127.84 via2_1600x480 ;
      VIA 264.1 127.84 via_1600x480 ;
      VIA 243.9 127.84 via3_1600x480 ;
      VIA 243.9 127.84 via2_1600x480 ;
      VIA 243.9 127.84 via_1600x480 ;
      VIA 223.7 127.84 via3_1600x480 ;
      VIA 223.7 127.84 via2_1600x480 ;
      VIA 223.7 127.84 via_1600x480 ;
      VIA 203.5 127.84 via3_1600x480 ;
      VIA 203.5 127.84 via2_1600x480 ;
      VIA 203.5 127.84 via_1600x480 ;
      VIA 183.3 127.84 via3_1600x480 ;
      VIA 183.3 127.84 via2_1600x480 ;
      VIA 183.3 127.84 via_1600x480 ;
      VIA 163.1 127.84 via3_1600x480 ;
      VIA 163.1 127.84 via2_1600x480 ;
      VIA 163.1 127.84 via_1600x480 ;
      VIA 142.9 127.84 via3_1600x480 ;
      VIA 142.9 127.84 via2_1600x480 ;
      VIA 142.9 127.84 via_1600x480 ;
      VIA 122.7 127.84 via3_1600x480 ;
      VIA 122.7 127.84 via2_1600x480 ;
      VIA 122.7 127.84 via_1600x480 ;
      VIA 102.5 127.84 via3_1600x480 ;
      VIA 102.5 127.84 via2_1600x480 ;
      VIA 102.5 127.84 via_1600x480 ;
      VIA 82.3 127.84 via3_1600x480 ;
      VIA 82.3 127.84 via2_1600x480 ;
      VIA 82.3 127.84 via_1600x480 ;
      VIA 62.1 127.84 via3_1600x480 ;
      VIA 62.1 127.84 via2_1600x480 ;
      VIA 62.1 127.84 via_1600x480 ;
      VIA 41.9 127.84 via3_1600x480 ;
      VIA 41.9 127.84 via2_1600x480 ;
      VIA 41.9 127.84 via_1600x480 ;
      VIA 21.7 127.84 via3_1600x480 ;
      VIA 21.7 127.84 via2_1600x480 ;
      VIA 21.7 127.84 via_1600x480 ;
      VIA 344.9 122.4 via3_1600x480 ;
      VIA 344.9 122.4 via2_1600x480 ;
      VIA 344.9 122.4 via_1600x480 ;
      VIA 324.7 122.4 via3_1600x480 ;
      VIA 324.7 122.4 via2_1600x480 ;
      VIA 324.7 122.4 via_1600x480 ;
      VIA 304.5 122.4 via3_1600x480 ;
      VIA 304.5 122.4 via2_1600x480 ;
      VIA 304.5 122.4 via_1600x480 ;
      VIA 284.3 122.4 via3_1600x480 ;
      VIA 284.3 122.4 via2_1600x480 ;
      VIA 284.3 122.4 via_1600x480 ;
      VIA 264.1 122.4 via3_1600x480 ;
      VIA 264.1 122.4 via2_1600x480 ;
      VIA 264.1 122.4 via_1600x480 ;
      VIA 243.9 122.4 via3_1600x480 ;
      VIA 243.9 122.4 via2_1600x480 ;
      VIA 243.9 122.4 via_1600x480 ;
      VIA 223.7 122.4 via3_1600x480 ;
      VIA 223.7 122.4 via2_1600x480 ;
      VIA 223.7 122.4 via_1600x480 ;
      VIA 203.5 122.4 via3_1600x480 ;
      VIA 203.5 122.4 via2_1600x480 ;
      VIA 203.5 122.4 via_1600x480 ;
      VIA 183.3 122.4 via3_1600x480 ;
      VIA 183.3 122.4 via2_1600x480 ;
      VIA 183.3 122.4 via_1600x480 ;
      VIA 163.1 122.4 via3_1600x480 ;
      VIA 163.1 122.4 via2_1600x480 ;
      VIA 163.1 122.4 via_1600x480 ;
      VIA 142.9 122.4 via3_1600x480 ;
      VIA 142.9 122.4 via2_1600x480 ;
      VIA 142.9 122.4 via_1600x480 ;
      VIA 122.7 122.4 via3_1600x480 ;
      VIA 122.7 122.4 via2_1600x480 ;
      VIA 122.7 122.4 via_1600x480 ;
      VIA 102.5 122.4 via3_1600x480 ;
      VIA 102.5 122.4 via2_1600x480 ;
      VIA 102.5 122.4 via_1600x480 ;
      VIA 82.3 122.4 via3_1600x480 ;
      VIA 82.3 122.4 via2_1600x480 ;
      VIA 82.3 122.4 via_1600x480 ;
      VIA 62.1 122.4 via3_1600x480 ;
      VIA 62.1 122.4 via2_1600x480 ;
      VIA 62.1 122.4 via_1600x480 ;
      VIA 41.9 122.4 via3_1600x480 ;
      VIA 41.9 122.4 via2_1600x480 ;
      VIA 41.9 122.4 via_1600x480 ;
      VIA 21.7 122.4 via3_1600x480 ;
      VIA 21.7 122.4 via2_1600x480 ;
      VIA 21.7 122.4 via_1600x480 ;
      VIA 344.9 116.96 via3_1600x480 ;
      VIA 344.9 116.96 via2_1600x480 ;
      VIA 344.9 116.96 via_1600x480 ;
      VIA 324.7 116.96 via3_1600x480 ;
      VIA 324.7 116.96 via2_1600x480 ;
      VIA 324.7 116.96 via_1600x480 ;
      VIA 304.5 116.96 via3_1600x480 ;
      VIA 304.5 116.96 via2_1600x480 ;
      VIA 304.5 116.96 via_1600x480 ;
      VIA 284.3 116.96 via3_1600x480 ;
      VIA 284.3 116.96 via2_1600x480 ;
      VIA 284.3 116.96 via_1600x480 ;
      VIA 264.1 116.96 via3_1600x480 ;
      VIA 264.1 116.96 via2_1600x480 ;
      VIA 264.1 116.96 via_1600x480 ;
      VIA 243.9 116.96 via3_1600x480 ;
      VIA 243.9 116.96 via2_1600x480 ;
      VIA 243.9 116.96 via_1600x480 ;
      VIA 223.7 116.96 via3_1600x480 ;
      VIA 223.7 116.96 via2_1600x480 ;
      VIA 223.7 116.96 via_1600x480 ;
      VIA 203.5 116.96 via3_1600x480 ;
      VIA 203.5 116.96 via2_1600x480 ;
      VIA 203.5 116.96 via_1600x480 ;
      VIA 183.3 116.96 via3_1600x480 ;
      VIA 183.3 116.96 via2_1600x480 ;
      VIA 183.3 116.96 via_1600x480 ;
      VIA 163.1 116.96 via3_1600x480 ;
      VIA 163.1 116.96 via2_1600x480 ;
      VIA 163.1 116.96 via_1600x480 ;
      VIA 142.9 116.96 via3_1600x480 ;
      VIA 142.9 116.96 via2_1600x480 ;
      VIA 142.9 116.96 via_1600x480 ;
      VIA 122.7 116.96 via3_1600x480 ;
      VIA 122.7 116.96 via2_1600x480 ;
      VIA 122.7 116.96 via_1600x480 ;
      VIA 102.5 116.96 via3_1600x480 ;
      VIA 102.5 116.96 via2_1600x480 ;
      VIA 102.5 116.96 via_1600x480 ;
      VIA 82.3 116.96 via3_1600x480 ;
      VIA 82.3 116.96 via2_1600x480 ;
      VIA 82.3 116.96 via_1600x480 ;
      VIA 62.1 116.96 via3_1600x480 ;
      VIA 62.1 116.96 via2_1600x480 ;
      VIA 62.1 116.96 via_1600x480 ;
      VIA 41.9 116.96 via3_1600x480 ;
      VIA 41.9 116.96 via2_1600x480 ;
      VIA 41.9 116.96 via_1600x480 ;
      VIA 21.7 116.96 via3_1600x480 ;
      VIA 21.7 116.96 via2_1600x480 ;
      VIA 21.7 116.96 via_1600x480 ;
      VIA 344.9 111.52 via3_1600x480 ;
      VIA 344.9 111.52 via2_1600x480 ;
      VIA 344.9 111.52 via_1600x480 ;
      VIA 324.7 111.52 via3_1600x480 ;
      VIA 324.7 111.52 via2_1600x480 ;
      VIA 324.7 111.52 via_1600x480 ;
      VIA 304.5 111.52 via3_1600x480 ;
      VIA 304.5 111.52 via2_1600x480 ;
      VIA 304.5 111.52 via_1600x480 ;
      VIA 284.3 111.52 via3_1600x480 ;
      VIA 284.3 111.52 via2_1600x480 ;
      VIA 284.3 111.52 via_1600x480 ;
      VIA 264.1 111.52 via3_1600x480 ;
      VIA 264.1 111.52 via2_1600x480 ;
      VIA 264.1 111.52 via_1600x480 ;
      VIA 243.9 111.52 via3_1600x480 ;
      VIA 243.9 111.52 via2_1600x480 ;
      VIA 243.9 111.52 via_1600x480 ;
      VIA 223.7 111.52 via3_1600x480 ;
      VIA 223.7 111.52 via2_1600x480 ;
      VIA 223.7 111.52 via_1600x480 ;
      VIA 203.5 111.52 via3_1600x480 ;
      VIA 203.5 111.52 via2_1600x480 ;
      VIA 203.5 111.52 via_1600x480 ;
      VIA 183.3 111.52 via3_1600x480 ;
      VIA 183.3 111.52 via2_1600x480 ;
      VIA 183.3 111.52 via_1600x480 ;
      VIA 163.1 111.52 via3_1600x480 ;
      VIA 163.1 111.52 via2_1600x480 ;
      VIA 163.1 111.52 via_1600x480 ;
      VIA 142.9 111.52 via3_1600x480 ;
      VIA 142.9 111.52 via2_1600x480 ;
      VIA 142.9 111.52 via_1600x480 ;
      VIA 122.7 111.52 via3_1600x480 ;
      VIA 122.7 111.52 via2_1600x480 ;
      VIA 122.7 111.52 via_1600x480 ;
      VIA 102.5 111.52 via3_1600x480 ;
      VIA 102.5 111.52 via2_1600x480 ;
      VIA 102.5 111.52 via_1600x480 ;
      VIA 82.3 111.52 via3_1600x480 ;
      VIA 82.3 111.52 via2_1600x480 ;
      VIA 82.3 111.52 via_1600x480 ;
      VIA 62.1 111.52 via3_1600x480 ;
      VIA 62.1 111.52 via2_1600x480 ;
      VIA 62.1 111.52 via_1600x480 ;
      VIA 41.9 111.52 via3_1600x480 ;
      VIA 41.9 111.52 via2_1600x480 ;
      VIA 41.9 111.52 via_1600x480 ;
      VIA 21.7 111.52 via3_1600x480 ;
      VIA 21.7 111.52 via2_1600x480 ;
      VIA 21.7 111.52 via_1600x480 ;
      VIA 344.9 106.08 via3_1600x480 ;
      VIA 344.9 106.08 via2_1600x480 ;
      VIA 344.9 106.08 via_1600x480 ;
      VIA 324.7 106.08 via3_1600x480 ;
      VIA 324.7 106.08 via2_1600x480 ;
      VIA 324.7 106.08 via_1600x480 ;
      VIA 304.5 106.08 via3_1600x480 ;
      VIA 304.5 106.08 via2_1600x480 ;
      VIA 304.5 106.08 via_1600x480 ;
      VIA 284.3 106.08 via3_1600x480 ;
      VIA 284.3 106.08 via2_1600x480 ;
      VIA 284.3 106.08 via_1600x480 ;
      VIA 264.1 106.08 via3_1600x480 ;
      VIA 264.1 106.08 via2_1600x480 ;
      VIA 264.1 106.08 via_1600x480 ;
      VIA 243.9 106.08 via3_1600x480 ;
      VIA 243.9 106.08 via2_1600x480 ;
      VIA 243.9 106.08 via_1600x480 ;
      VIA 223.7 106.08 via3_1600x480 ;
      VIA 223.7 106.08 via2_1600x480 ;
      VIA 223.7 106.08 via_1600x480 ;
      VIA 203.5 106.08 via3_1600x480 ;
      VIA 203.5 106.08 via2_1600x480 ;
      VIA 203.5 106.08 via_1600x480 ;
      VIA 183.3 106.08 via3_1600x480 ;
      VIA 183.3 106.08 via2_1600x480 ;
      VIA 183.3 106.08 via_1600x480 ;
      VIA 163.1 106.08 via3_1600x480 ;
      VIA 163.1 106.08 via2_1600x480 ;
      VIA 163.1 106.08 via_1600x480 ;
      VIA 142.9 106.08 via3_1600x480 ;
      VIA 142.9 106.08 via2_1600x480 ;
      VIA 142.9 106.08 via_1600x480 ;
      VIA 122.7 106.08 via3_1600x480 ;
      VIA 122.7 106.08 via2_1600x480 ;
      VIA 122.7 106.08 via_1600x480 ;
      VIA 102.5 106.08 via3_1600x480 ;
      VIA 102.5 106.08 via2_1600x480 ;
      VIA 102.5 106.08 via_1600x480 ;
      VIA 82.3 106.08 via3_1600x480 ;
      VIA 82.3 106.08 via2_1600x480 ;
      VIA 82.3 106.08 via_1600x480 ;
      VIA 62.1 106.08 via3_1600x480 ;
      VIA 62.1 106.08 via2_1600x480 ;
      VIA 62.1 106.08 via_1600x480 ;
      VIA 41.9 106.08 via3_1600x480 ;
      VIA 41.9 106.08 via2_1600x480 ;
      VIA 41.9 106.08 via_1600x480 ;
      VIA 21.7 106.08 via3_1600x480 ;
      VIA 21.7 106.08 via2_1600x480 ;
      VIA 21.7 106.08 via_1600x480 ;
      VIA 344.9 100.64 via3_1600x480 ;
      VIA 344.9 100.64 via2_1600x480 ;
      VIA 344.9 100.64 via_1600x480 ;
      VIA 324.7 100.64 via3_1600x480 ;
      VIA 324.7 100.64 via2_1600x480 ;
      VIA 324.7 100.64 via_1600x480 ;
      VIA 304.5 100.64 via3_1600x480 ;
      VIA 304.5 100.64 via2_1600x480 ;
      VIA 304.5 100.64 via_1600x480 ;
      VIA 284.3 100.64 via3_1600x480 ;
      VIA 284.3 100.64 via2_1600x480 ;
      VIA 284.3 100.64 via_1600x480 ;
      VIA 264.1 100.64 via3_1600x480 ;
      VIA 264.1 100.64 via2_1600x480 ;
      VIA 264.1 100.64 via_1600x480 ;
      VIA 243.9 100.64 via3_1600x480 ;
      VIA 243.9 100.64 via2_1600x480 ;
      VIA 243.9 100.64 via_1600x480 ;
      VIA 223.7 100.64 via3_1600x480 ;
      VIA 223.7 100.64 via2_1600x480 ;
      VIA 223.7 100.64 via_1600x480 ;
      VIA 203.5 100.64 via3_1600x480 ;
      VIA 203.5 100.64 via2_1600x480 ;
      VIA 203.5 100.64 via_1600x480 ;
      VIA 183.3 100.64 via3_1600x480 ;
      VIA 183.3 100.64 via2_1600x480 ;
      VIA 183.3 100.64 via_1600x480 ;
      VIA 163.1 100.64 via3_1600x480 ;
      VIA 163.1 100.64 via2_1600x480 ;
      VIA 163.1 100.64 via_1600x480 ;
      VIA 142.9 100.64 via3_1600x480 ;
      VIA 142.9 100.64 via2_1600x480 ;
      VIA 142.9 100.64 via_1600x480 ;
      VIA 122.7 100.64 via3_1600x480 ;
      VIA 122.7 100.64 via2_1600x480 ;
      VIA 122.7 100.64 via_1600x480 ;
      VIA 102.5 100.64 via3_1600x480 ;
      VIA 102.5 100.64 via2_1600x480 ;
      VIA 102.5 100.64 via_1600x480 ;
      VIA 82.3 100.64 via3_1600x480 ;
      VIA 82.3 100.64 via2_1600x480 ;
      VIA 82.3 100.64 via_1600x480 ;
      VIA 62.1 100.64 via3_1600x480 ;
      VIA 62.1 100.64 via2_1600x480 ;
      VIA 62.1 100.64 via_1600x480 ;
      VIA 41.9 100.64 via3_1600x480 ;
      VIA 41.9 100.64 via2_1600x480 ;
      VIA 41.9 100.64 via_1600x480 ;
      VIA 21.7 100.64 via3_1600x480 ;
      VIA 21.7 100.64 via2_1600x480 ;
      VIA 21.7 100.64 via_1600x480 ;
      VIA 344.9 95.2 via3_1600x480 ;
      VIA 344.9 95.2 via2_1600x480 ;
      VIA 344.9 95.2 via_1600x480 ;
      VIA 324.7 95.2 via3_1600x480 ;
      VIA 324.7 95.2 via2_1600x480 ;
      VIA 324.7 95.2 via_1600x480 ;
      VIA 304.5 95.2 via3_1600x480 ;
      VIA 304.5 95.2 via2_1600x480 ;
      VIA 304.5 95.2 via_1600x480 ;
      VIA 284.3 95.2 via3_1600x480 ;
      VIA 284.3 95.2 via2_1600x480 ;
      VIA 284.3 95.2 via_1600x480 ;
      VIA 264.1 95.2 via3_1600x480 ;
      VIA 264.1 95.2 via2_1600x480 ;
      VIA 264.1 95.2 via_1600x480 ;
      VIA 243.9 95.2 via3_1600x480 ;
      VIA 243.9 95.2 via2_1600x480 ;
      VIA 243.9 95.2 via_1600x480 ;
      VIA 223.7 95.2 via3_1600x480 ;
      VIA 223.7 95.2 via2_1600x480 ;
      VIA 223.7 95.2 via_1600x480 ;
      VIA 203.5 95.2 via3_1600x480 ;
      VIA 203.5 95.2 via2_1600x480 ;
      VIA 203.5 95.2 via_1600x480 ;
      VIA 183.3 95.2 via3_1600x480 ;
      VIA 183.3 95.2 via2_1600x480 ;
      VIA 183.3 95.2 via_1600x480 ;
      VIA 163.1 95.2 via3_1600x480 ;
      VIA 163.1 95.2 via2_1600x480 ;
      VIA 163.1 95.2 via_1600x480 ;
      VIA 142.9 95.2 via3_1600x480 ;
      VIA 142.9 95.2 via2_1600x480 ;
      VIA 142.9 95.2 via_1600x480 ;
      VIA 122.7 95.2 via3_1600x480 ;
      VIA 122.7 95.2 via2_1600x480 ;
      VIA 122.7 95.2 via_1600x480 ;
      VIA 102.5 95.2 via3_1600x480 ;
      VIA 102.5 95.2 via2_1600x480 ;
      VIA 102.5 95.2 via_1600x480 ;
      VIA 82.3 95.2 via3_1600x480 ;
      VIA 82.3 95.2 via2_1600x480 ;
      VIA 82.3 95.2 via_1600x480 ;
      VIA 62.1 95.2 via3_1600x480 ;
      VIA 62.1 95.2 via2_1600x480 ;
      VIA 62.1 95.2 via_1600x480 ;
      VIA 41.9 95.2 via3_1600x480 ;
      VIA 41.9 95.2 via2_1600x480 ;
      VIA 41.9 95.2 via_1600x480 ;
      VIA 21.7 95.2 via3_1600x480 ;
      VIA 21.7 95.2 via2_1600x480 ;
      VIA 21.7 95.2 via_1600x480 ;
      VIA 344.9 89.76 via3_1600x480 ;
      VIA 344.9 89.76 via2_1600x480 ;
      VIA 344.9 89.76 via_1600x480 ;
      VIA 324.7 89.76 via3_1600x480 ;
      VIA 324.7 89.76 via2_1600x480 ;
      VIA 324.7 89.76 via_1600x480 ;
      VIA 304.5 89.76 via3_1600x480 ;
      VIA 304.5 89.76 via2_1600x480 ;
      VIA 304.5 89.76 via_1600x480 ;
      VIA 284.3 89.76 via3_1600x480 ;
      VIA 284.3 89.76 via2_1600x480 ;
      VIA 284.3 89.76 via_1600x480 ;
      VIA 264.1 89.76 via3_1600x480 ;
      VIA 264.1 89.76 via2_1600x480 ;
      VIA 264.1 89.76 via_1600x480 ;
      VIA 243.9 89.76 via3_1600x480 ;
      VIA 243.9 89.76 via2_1600x480 ;
      VIA 243.9 89.76 via_1600x480 ;
      VIA 223.7 89.76 via3_1600x480 ;
      VIA 223.7 89.76 via2_1600x480 ;
      VIA 223.7 89.76 via_1600x480 ;
      VIA 203.5 89.76 via3_1600x480 ;
      VIA 203.5 89.76 via2_1600x480 ;
      VIA 203.5 89.76 via_1600x480 ;
      VIA 183.3 89.76 via3_1600x480 ;
      VIA 183.3 89.76 via2_1600x480 ;
      VIA 183.3 89.76 via_1600x480 ;
      VIA 163.1 89.76 via3_1600x480 ;
      VIA 163.1 89.76 via2_1600x480 ;
      VIA 163.1 89.76 via_1600x480 ;
      VIA 142.9 89.76 via3_1600x480 ;
      VIA 142.9 89.76 via2_1600x480 ;
      VIA 142.9 89.76 via_1600x480 ;
      VIA 122.7 89.76 via3_1600x480 ;
      VIA 122.7 89.76 via2_1600x480 ;
      VIA 122.7 89.76 via_1600x480 ;
      VIA 102.5 89.76 via3_1600x480 ;
      VIA 102.5 89.76 via2_1600x480 ;
      VIA 102.5 89.76 via_1600x480 ;
      VIA 82.3 89.76 via3_1600x480 ;
      VIA 82.3 89.76 via2_1600x480 ;
      VIA 82.3 89.76 via_1600x480 ;
      VIA 62.1 89.76 via3_1600x480 ;
      VIA 62.1 89.76 via2_1600x480 ;
      VIA 62.1 89.76 via_1600x480 ;
      VIA 41.9 89.76 via3_1600x480 ;
      VIA 41.9 89.76 via2_1600x480 ;
      VIA 41.9 89.76 via_1600x480 ;
      VIA 21.7 89.76 via3_1600x480 ;
      VIA 21.7 89.76 via2_1600x480 ;
      VIA 21.7 89.76 via_1600x480 ;
      VIA 344.9 84.32 via3_1600x480 ;
      VIA 344.9 84.32 via2_1600x480 ;
      VIA 344.9 84.32 via_1600x480 ;
      VIA 324.7 84.32 via3_1600x480 ;
      VIA 324.7 84.32 via2_1600x480 ;
      VIA 324.7 84.32 via_1600x480 ;
      VIA 304.5 84.32 via3_1600x480 ;
      VIA 304.5 84.32 via2_1600x480 ;
      VIA 304.5 84.32 via_1600x480 ;
      VIA 284.3 84.32 via3_1600x480 ;
      VIA 284.3 84.32 via2_1600x480 ;
      VIA 284.3 84.32 via_1600x480 ;
      VIA 264.1 84.32 via3_1600x480 ;
      VIA 264.1 84.32 via2_1600x480 ;
      VIA 264.1 84.32 via_1600x480 ;
      VIA 243.9 84.32 via3_1600x480 ;
      VIA 243.9 84.32 via2_1600x480 ;
      VIA 243.9 84.32 via_1600x480 ;
      VIA 223.7 84.32 via3_1600x480 ;
      VIA 223.7 84.32 via2_1600x480 ;
      VIA 223.7 84.32 via_1600x480 ;
      VIA 203.5 84.32 via3_1600x480 ;
      VIA 203.5 84.32 via2_1600x480 ;
      VIA 203.5 84.32 via_1600x480 ;
      VIA 183.3 84.32 via3_1600x480 ;
      VIA 183.3 84.32 via2_1600x480 ;
      VIA 183.3 84.32 via_1600x480 ;
      VIA 163.1 84.32 via3_1600x480 ;
      VIA 163.1 84.32 via2_1600x480 ;
      VIA 163.1 84.32 via_1600x480 ;
      VIA 142.9 84.32 via3_1600x480 ;
      VIA 142.9 84.32 via2_1600x480 ;
      VIA 142.9 84.32 via_1600x480 ;
      VIA 122.7 84.32 via3_1600x480 ;
      VIA 122.7 84.32 via2_1600x480 ;
      VIA 122.7 84.32 via_1600x480 ;
      VIA 102.5 84.32 via3_1600x480 ;
      VIA 102.5 84.32 via2_1600x480 ;
      VIA 102.5 84.32 via_1600x480 ;
      VIA 82.3 84.32 via3_1600x480 ;
      VIA 82.3 84.32 via2_1600x480 ;
      VIA 82.3 84.32 via_1600x480 ;
      VIA 62.1 84.32 via3_1600x480 ;
      VIA 62.1 84.32 via2_1600x480 ;
      VIA 62.1 84.32 via_1600x480 ;
      VIA 41.9 84.32 via3_1600x480 ;
      VIA 41.9 84.32 via2_1600x480 ;
      VIA 41.9 84.32 via_1600x480 ;
      VIA 21.7 84.32 via3_1600x480 ;
      VIA 21.7 84.32 via2_1600x480 ;
      VIA 21.7 84.32 via_1600x480 ;
      VIA 344.9 78.88 via3_1600x480 ;
      VIA 344.9 78.88 via2_1600x480 ;
      VIA 344.9 78.88 via_1600x480 ;
      VIA 324.7 78.88 via3_1600x480 ;
      VIA 324.7 78.88 via2_1600x480 ;
      VIA 324.7 78.88 via_1600x480 ;
      VIA 304.5 78.88 via3_1600x480 ;
      VIA 304.5 78.88 via2_1600x480 ;
      VIA 304.5 78.88 via_1600x480 ;
      VIA 284.3 78.88 via3_1600x480 ;
      VIA 284.3 78.88 via2_1600x480 ;
      VIA 284.3 78.88 via_1600x480 ;
      VIA 264.1 78.88 via3_1600x480 ;
      VIA 264.1 78.88 via2_1600x480 ;
      VIA 264.1 78.88 via_1600x480 ;
      VIA 243.9 78.88 via3_1600x480 ;
      VIA 243.9 78.88 via2_1600x480 ;
      VIA 243.9 78.88 via_1600x480 ;
      VIA 223.7 78.88 via3_1600x480 ;
      VIA 223.7 78.88 via2_1600x480 ;
      VIA 223.7 78.88 via_1600x480 ;
      VIA 203.5 78.88 via3_1600x480 ;
      VIA 203.5 78.88 via2_1600x480 ;
      VIA 203.5 78.88 via_1600x480 ;
      VIA 183.3 78.88 via3_1600x480 ;
      VIA 183.3 78.88 via2_1600x480 ;
      VIA 183.3 78.88 via_1600x480 ;
      VIA 163.1 78.88 via3_1600x480 ;
      VIA 163.1 78.88 via2_1600x480 ;
      VIA 163.1 78.88 via_1600x480 ;
      VIA 142.9 78.88 via3_1600x480 ;
      VIA 142.9 78.88 via2_1600x480 ;
      VIA 142.9 78.88 via_1600x480 ;
      VIA 122.7 78.88 via3_1600x480 ;
      VIA 122.7 78.88 via2_1600x480 ;
      VIA 122.7 78.88 via_1600x480 ;
      VIA 102.5 78.88 via3_1600x480 ;
      VIA 102.5 78.88 via2_1600x480 ;
      VIA 102.5 78.88 via_1600x480 ;
      VIA 82.3 78.88 via3_1600x480 ;
      VIA 82.3 78.88 via2_1600x480 ;
      VIA 82.3 78.88 via_1600x480 ;
      VIA 62.1 78.88 via3_1600x480 ;
      VIA 62.1 78.88 via2_1600x480 ;
      VIA 62.1 78.88 via_1600x480 ;
      VIA 41.9 78.88 via3_1600x480 ;
      VIA 41.9 78.88 via2_1600x480 ;
      VIA 41.9 78.88 via_1600x480 ;
      VIA 21.7 78.88 via3_1600x480 ;
      VIA 21.7 78.88 via2_1600x480 ;
      VIA 21.7 78.88 via_1600x480 ;
      VIA 344.9 73.44 via3_1600x480 ;
      VIA 344.9 73.44 via2_1600x480 ;
      VIA 344.9 73.44 via_1600x480 ;
      VIA 324.7 73.44 via3_1600x480 ;
      VIA 324.7 73.44 via2_1600x480 ;
      VIA 324.7 73.44 via_1600x480 ;
      VIA 304.5 73.44 via3_1600x480 ;
      VIA 304.5 73.44 via2_1600x480 ;
      VIA 304.5 73.44 via_1600x480 ;
      VIA 284.3 73.44 via3_1600x480 ;
      VIA 284.3 73.44 via2_1600x480 ;
      VIA 284.3 73.44 via_1600x480 ;
      VIA 264.1 73.44 via3_1600x480 ;
      VIA 264.1 73.44 via2_1600x480 ;
      VIA 264.1 73.44 via_1600x480 ;
      VIA 243.9 73.44 via3_1600x480 ;
      VIA 243.9 73.44 via2_1600x480 ;
      VIA 243.9 73.44 via_1600x480 ;
      VIA 223.7 73.44 via3_1600x480 ;
      VIA 223.7 73.44 via2_1600x480 ;
      VIA 223.7 73.44 via_1600x480 ;
      VIA 203.5 73.44 via3_1600x480 ;
      VIA 203.5 73.44 via2_1600x480 ;
      VIA 203.5 73.44 via_1600x480 ;
      VIA 183.3 73.44 via3_1600x480 ;
      VIA 183.3 73.44 via2_1600x480 ;
      VIA 183.3 73.44 via_1600x480 ;
      VIA 163.1 73.44 via3_1600x480 ;
      VIA 163.1 73.44 via2_1600x480 ;
      VIA 163.1 73.44 via_1600x480 ;
      VIA 142.9 73.44 via3_1600x480 ;
      VIA 142.9 73.44 via2_1600x480 ;
      VIA 142.9 73.44 via_1600x480 ;
      VIA 122.7 73.44 via3_1600x480 ;
      VIA 122.7 73.44 via2_1600x480 ;
      VIA 122.7 73.44 via_1600x480 ;
      VIA 102.5 73.44 via3_1600x480 ;
      VIA 102.5 73.44 via2_1600x480 ;
      VIA 102.5 73.44 via_1600x480 ;
      VIA 82.3 73.44 via3_1600x480 ;
      VIA 82.3 73.44 via2_1600x480 ;
      VIA 82.3 73.44 via_1600x480 ;
      VIA 62.1 73.44 via3_1600x480 ;
      VIA 62.1 73.44 via2_1600x480 ;
      VIA 62.1 73.44 via_1600x480 ;
      VIA 41.9 73.44 via3_1600x480 ;
      VIA 41.9 73.44 via2_1600x480 ;
      VIA 41.9 73.44 via_1600x480 ;
      VIA 21.7 73.44 via3_1600x480 ;
      VIA 21.7 73.44 via2_1600x480 ;
      VIA 21.7 73.44 via_1600x480 ;
      VIA 344.9 68 via3_1600x480 ;
      VIA 344.9 68 via2_1600x480 ;
      VIA 344.9 68 via_1600x480 ;
      VIA 324.7 68 via3_1600x480 ;
      VIA 324.7 68 via2_1600x480 ;
      VIA 324.7 68 via_1600x480 ;
      VIA 304.5 68 via3_1600x480 ;
      VIA 304.5 68 via2_1600x480 ;
      VIA 304.5 68 via_1600x480 ;
      VIA 284.3 68 via3_1600x480 ;
      VIA 284.3 68 via2_1600x480 ;
      VIA 284.3 68 via_1600x480 ;
      VIA 264.1 68 via3_1600x480 ;
      VIA 264.1 68 via2_1600x480 ;
      VIA 264.1 68 via_1600x480 ;
      VIA 243.9 68 via3_1600x480 ;
      VIA 243.9 68 via2_1600x480 ;
      VIA 243.9 68 via_1600x480 ;
      VIA 223.7 68 via3_1600x480 ;
      VIA 223.7 68 via2_1600x480 ;
      VIA 223.7 68 via_1600x480 ;
      VIA 203.5 68 via3_1600x480 ;
      VIA 203.5 68 via2_1600x480 ;
      VIA 203.5 68 via_1600x480 ;
      VIA 183.3 68 via3_1600x480 ;
      VIA 183.3 68 via2_1600x480 ;
      VIA 183.3 68 via_1600x480 ;
      VIA 163.1 68 via3_1600x480 ;
      VIA 163.1 68 via2_1600x480 ;
      VIA 163.1 68 via_1600x480 ;
      VIA 142.9 68 via3_1600x480 ;
      VIA 142.9 68 via2_1600x480 ;
      VIA 142.9 68 via_1600x480 ;
      VIA 122.7 68 via3_1600x480 ;
      VIA 122.7 68 via2_1600x480 ;
      VIA 122.7 68 via_1600x480 ;
      VIA 102.5 68 via3_1600x480 ;
      VIA 102.5 68 via2_1600x480 ;
      VIA 102.5 68 via_1600x480 ;
      VIA 82.3 68 via3_1600x480 ;
      VIA 82.3 68 via2_1600x480 ;
      VIA 82.3 68 via_1600x480 ;
      VIA 62.1 68 via3_1600x480 ;
      VIA 62.1 68 via2_1600x480 ;
      VIA 62.1 68 via_1600x480 ;
      VIA 41.9 68 via3_1600x480 ;
      VIA 41.9 68 via2_1600x480 ;
      VIA 41.9 68 via_1600x480 ;
      VIA 21.7 68 via3_1600x480 ;
      VIA 21.7 68 via2_1600x480 ;
      VIA 21.7 68 via_1600x480 ;
      VIA 344.9 62.56 via3_1600x480 ;
      VIA 344.9 62.56 via2_1600x480 ;
      VIA 344.9 62.56 via_1600x480 ;
      VIA 324.7 62.56 via3_1600x480 ;
      VIA 324.7 62.56 via2_1600x480 ;
      VIA 324.7 62.56 via_1600x480 ;
      VIA 304.5 62.56 via3_1600x480 ;
      VIA 304.5 62.56 via2_1600x480 ;
      VIA 304.5 62.56 via_1600x480 ;
      VIA 284.3 62.56 via3_1600x480 ;
      VIA 284.3 62.56 via2_1600x480 ;
      VIA 284.3 62.56 via_1600x480 ;
      VIA 264.1 62.56 via3_1600x480 ;
      VIA 264.1 62.56 via2_1600x480 ;
      VIA 264.1 62.56 via_1600x480 ;
      VIA 243.9 62.56 via3_1600x480 ;
      VIA 243.9 62.56 via2_1600x480 ;
      VIA 243.9 62.56 via_1600x480 ;
      VIA 223.7 62.56 via3_1600x480 ;
      VIA 223.7 62.56 via2_1600x480 ;
      VIA 223.7 62.56 via_1600x480 ;
      VIA 203.5 62.56 via3_1600x480 ;
      VIA 203.5 62.56 via2_1600x480 ;
      VIA 203.5 62.56 via_1600x480 ;
      VIA 183.3 62.56 via3_1600x480 ;
      VIA 183.3 62.56 via2_1600x480 ;
      VIA 183.3 62.56 via_1600x480 ;
      VIA 163.1 62.56 via3_1600x480 ;
      VIA 163.1 62.56 via2_1600x480 ;
      VIA 163.1 62.56 via_1600x480 ;
      VIA 142.9 62.56 via3_1600x480 ;
      VIA 142.9 62.56 via2_1600x480 ;
      VIA 142.9 62.56 via_1600x480 ;
      VIA 122.7 62.56 via3_1600x480 ;
      VIA 122.7 62.56 via2_1600x480 ;
      VIA 122.7 62.56 via_1600x480 ;
      VIA 102.5 62.56 via3_1600x480 ;
      VIA 102.5 62.56 via2_1600x480 ;
      VIA 102.5 62.56 via_1600x480 ;
      VIA 82.3 62.56 via3_1600x480 ;
      VIA 82.3 62.56 via2_1600x480 ;
      VIA 82.3 62.56 via_1600x480 ;
      VIA 62.1 62.56 via3_1600x480 ;
      VIA 62.1 62.56 via2_1600x480 ;
      VIA 62.1 62.56 via_1600x480 ;
      VIA 41.9 62.56 via3_1600x480 ;
      VIA 41.9 62.56 via2_1600x480 ;
      VIA 41.9 62.56 via_1600x480 ;
      VIA 21.7 62.56 via3_1600x480 ;
      VIA 21.7 62.56 via2_1600x480 ;
      VIA 21.7 62.56 via_1600x480 ;
      VIA 344.9 57.12 via3_1600x480 ;
      VIA 344.9 57.12 via2_1600x480 ;
      VIA 344.9 57.12 via_1600x480 ;
      VIA 324.7 57.12 via3_1600x480 ;
      VIA 324.7 57.12 via2_1600x480 ;
      VIA 324.7 57.12 via_1600x480 ;
      VIA 304.5 57.12 via3_1600x480 ;
      VIA 304.5 57.12 via2_1600x480 ;
      VIA 304.5 57.12 via_1600x480 ;
      VIA 284.3 57.12 via3_1600x480 ;
      VIA 284.3 57.12 via2_1600x480 ;
      VIA 284.3 57.12 via_1600x480 ;
      VIA 264.1 57.12 via3_1600x480 ;
      VIA 264.1 57.12 via2_1600x480 ;
      VIA 264.1 57.12 via_1600x480 ;
      VIA 243.9 57.12 via3_1600x480 ;
      VIA 243.9 57.12 via2_1600x480 ;
      VIA 243.9 57.12 via_1600x480 ;
      VIA 223.7 57.12 via3_1600x480 ;
      VIA 223.7 57.12 via2_1600x480 ;
      VIA 223.7 57.12 via_1600x480 ;
      VIA 203.5 57.12 via3_1600x480 ;
      VIA 203.5 57.12 via2_1600x480 ;
      VIA 203.5 57.12 via_1600x480 ;
      VIA 183.3 57.12 via3_1600x480 ;
      VIA 183.3 57.12 via2_1600x480 ;
      VIA 183.3 57.12 via_1600x480 ;
      VIA 163.1 57.12 via3_1600x480 ;
      VIA 163.1 57.12 via2_1600x480 ;
      VIA 163.1 57.12 via_1600x480 ;
      VIA 142.9 57.12 via3_1600x480 ;
      VIA 142.9 57.12 via2_1600x480 ;
      VIA 142.9 57.12 via_1600x480 ;
      VIA 122.7 57.12 via3_1600x480 ;
      VIA 122.7 57.12 via2_1600x480 ;
      VIA 122.7 57.12 via_1600x480 ;
      VIA 102.5 57.12 via3_1600x480 ;
      VIA 102.5 57.12 via2_1600x480 ;
      VIA 102.5 57.12 via_1600x480 ;
      VIA 82.3 57.12 via3_1600x480 ;
      VIA 82.3 57.12 via2_1600x480 ;
      VIA 82.3 57.12 via_1600x480 ;
      VIA 62.1 57.12 via3_1600x480 ;
      VIA 62.1 57.12 via2_1600x480 ;
      VIA 62.1 57.12 via_1600x480 ;
      VIA 41.9 57.12 via3_1600x480 ;
      VIA 41.9 57.12 via2_1600x480 ;
      VIA 41.9 57.12 via_1600x480 ;
      VIA 21.7 57.12 via3_1600x480 ;
      VIA 21.7 57.12 via2_1600x480 ;
      VIA 21.7 57.12 via_1600x480 ;
      VIA 344.9 51.68 via3_1600x480 ;
      VIA 344.9 51.68 via2_1600x480 ;
      VIA 344.9 51.68 via_1600x480 ;
      VIA 324.7 51.68 via3_1600x480 ;
      VIA 324.7 51.68 via2_1600x480 ;
      VIA 324.7 51.68 via_1600x480 ;
      VIA 304.5 51.68 via3_1600x480 ;
      VIA 304.5 51.68 via2_1600x480 ;
      VIA 304.5 51.68 via_1600x480 ;
      VIA 284.3 51.68 via3_1600x480 ;
      VIA 284.3 51.68 via2_1600x480 ;
      VIA 284.3 51.68 via_1600x480 ;
      VIA 264.1 51.68 via3_1600x480 ;
      VIA 264.1 51.68 via2_1600x480 ;
      VIA 264.1 51.68 via_1600x480 ;
      VIA 243.9 51.68 via3_1600x480 ;
      VIA 243.9 51.68 via2_1600x480 ;
      VIA 243.9 51.68 via_1600x480 ;
      VIA 223.7 51.68 via3_1600x480 ;
      VIA 223.7 51.68 via2_1600x480 ;
      VIA 223.7 51.68 via_1600x480 ;
      VIA 203.5 51.68 via3_1600x480 ;
      VIA 203.5 51.68 via2_1600x480 ;
      VIA 203.5 51.68 via_1600x480 ;
      VIA 183.3 51.68 via3_1600x480 ;
      VIA 183.3 51.68 via2_1600x480 ;
      VIA 183.3 51.68 via_1600x480 ;
      VIA 163.1 51.68 via3_1600x480 ;
      VIA 163.1 51.68 via2_1600x480 ;
      VIA 163.1 51.68 via_1600x480 ;
      VIA 142.9 51.68 via3_1600x480 ;
      VIA 142.9 51.68 via2_1600x480 ;
      VIA 142.9 51.68 via_1600x480 ;
      VIA 122.7 51.68 via3_1600x480 ;
      VIA 122.7 51.68 via2_1600x480 ;
      VIA 122.7 51.68 via_1600x480 ;
      VIA 102.5 51.68 via3_1600x480 ;
      VIA 102.5 51.68 via2_1600x480 ;
      VIA 102.5 51.68 via_1600x480 ;
      VIA 82.3 51.68 via3_1600x480 ;
      VIA 82.3 51.68 via2_1600x480 ;
      VIA 82.3 51.68 via_1600x480 ;
      VIA 62.1 51.68 via3_1600x480 ;
      VIA 62.1 51.68 via2_1600x480 ;
      VIA 62.1 51.68 via_1600x480 ;
      VIA 41.9 51.68 via3_1600x480 ;
      VIA 41.9 51.68 via2_1600x480 ;
      VIA 41.9 51.68 via_1600x480 ;
      VIA 21.7 51.68 via3_1600x480 ;
      VIA 21.7 51.68 via2_1600x480 ;
      VIA 21.7 51.68 via_1600x480 ;
      VIA 344.9 46.24 via3_1600x480 ;
      VIA 344.9 46.24 via2_1600x480 ;
      VIA 344.9 46.24 via_1600x480 ;
      VIA 324.7 46.24 via3_1600x480 ;
      VIA 324.7 46.24 via2_1600x480 ;
      VIA 324.7 46.24 via_1600x480 ;
      VIA 304.5 46.24 via3_1600x480 ;
      VIA 304.5 46.24 via2_1600x480 ;
      VIA 304.5 46.24 via_1600x480 ;
      VIA 284.3 46.24 via3_1600x480 ;
      VIA 284.3 46.24 via2_1600x480 ;
      VIA 284.3 46.24 via_1600x480 ;
      VIA 264.1 46.24 via3_1600x480 ;
      VIA 264.1 46.24 via2_1600x480 ;
      VIA 264.1 46.24 via_1600x480 ;
      VIA 243.9 46.24 via3_1600x480 ;
      VIA 243.9 46.24 via2_1600x480 ;
      VIA 243.9 46.24 via_1600x480 ;
      VIA 223.7 46.24 via3_1600x480 ;
      VIA 223.7 46.24 via2_1600x480 ;
      VIA 223.7 46.24 via_1600x480 ;
      VIA 203.5 46.24 via3_1600x480 ;
      VIA 203.5 46.24 via2_1600x480 ;
      VIA 203.5 46.24 via_1600x480 ;
      VIA 183.3 46.24 via3_1600x480 ;
      VIA 183.3 46.24 via2_1600x480 ;
      VIA 183.3 46.24 via_1600x480 ;
      VIA 163.1 46.24 via3_1600x480 ;
      VIA 163.1 46.24 via2_1600x480 ;
      VIA 163.1 46.24 via_1600x480 ;
      VIA 142.9 46.24 via3_1600x480 ;
      VIA 142.9 46.24 via2_1600x480 ;
      VIA 142.9 46.24 via_1600x480 ;
      VIA 122.7 46.24 via3_1600x480 ;
      VIA 122.7 46.24 via2_1600x480 ;
      VIA 122.7 46.24 via_1600x480 ;
      VIA 102.5 46.24 via3_1600x480 ;
      VIA 102.5 46.24 via2_1600x480 ;
      VIA 102.5 46.24 via_1600x480 ;
      VIA 82.3 46.24 via3_1600x480 ;
      VIA 82.3 46.24 via2_1600x480 ;
      VIA 82.3 46.24 via_1600x480 ;
      VIA 62.1 46.24 via3_1600x480 ;
      VIA 62.1 46.24 via2_1600x480 ;
      VIA 62.1 46.24 via_1600x480 ;
      VIA 41.9 46.24 via3_1600x480 ;
      VIA 41.9 46.24 via2_1600x480 ;
      VIA 41.9 46.24 via_1600x480 ;
      VIA 21.7 46.24 via3_1600x480 ;
      VIA 21.7 46.24 via2_1600x480 ;
      VIA 21.7 46.24 via_1600x480 ;
      VIA 344.9 40.8 via3_1600x480 ;
      VIA 344.9 40.8 via2_1600x480 ;
      VIA 344.9 40.8 via_1600x480 ;
      VIA 324.7 40.8 via3_1600x480 ;
      VIA 324.7 40.8 via2_1600x480 ;
      VIA 324.7 40.8 via_1600x480 ;
      VIA 304.5 40.8 via3_1600x480 ;
      VIA 304.5 40.8 via2_1600x480 ;
      VIA 304.5 40.8 via_1600x480 ;
      VIA 284.3 40.8 via3_1600x480 ;
      VIA 284.3 40.8 via2_1600x480 ;
      VIA 284.3 40.8 via_1600x480 ;
      VIA 264.1 40.8 via3_1600x480 ;
      VIA 264.1 40.8 via2_1600x480 ;
      VIA 264.1 40.8 via_1600x480 ;
      VIA 243.9 40.8 via3_1600x480 ;
      VIA 243.9 40.8 via2_1600x480 ;
      VIA 243.9 40.8 via_1600x480 ;
      VIA 223.7 40.8 via3_1600x480 ;
      VIA 223.7 40.8 via2_1600x480 ;
      VIA 223.7 40.8 via_1600x480 ;
      VIA 203.5 40.8 via3_1600x480 ;
      VIA 203.5 40.8 via2_1600x480 ;
      VIA 203.5 40.8 via_1600x480 ;
      VIA 183.3 40.8 via3_1600x480 ;
      VIA 183.3 40.8 via2_1600x480 ;
      VIA 183.3 40.8 via_1600x480 ;
      VIA 163.1 40.8 via3_1600x480 ;
      VIA 163.1 40.8 via2_1600x480 ;
      VIA 163.1 40.8 via_1600x480 ;
      VIA 142.9 40.8 via3_1600x480 ;
      VIA 142.9 40.8 via2_1600x480 ;
      VIA 142.9 40.8 via_1600x480 ;
      VIA 122.7 40.8 via3_1600x480 ;
      VIA 122.7 40.8 via2_1600x480 ;
      VIA 122.7 40.8 via_1600x480 ;
      VIA 102.5 40.8 via3_1600x480 ;
      VIA 102.5 40.8 via2_1600x480 ;
      VIA 102.5 40.8 via_1600x480 ;
      VIA 82.3 40.8 via3_1600x480 ;
      VIA 82.3 40.8 via2_1600x480 ;
      VIA 82.3 40.8 via_1600x480 ;
      VIA 62.1 40.8 via3_1600x480 ;
      VIA 62.1 40.8 via2_1600x480 ;
      VIA 62.1 40.8 via_1600x480 ;
      VIA 41.9 40.8 via3_1600x480 ;
      VIA 41.9 40.8 via2_1600x480 ;
      VIA 41.9 40.8 via_1600x480 ;
      VIA 21.7 40.8 via3_1600x480 ;
      VIA 21.7 40.8 via2_1600x480 ;
      VIA 21.7 40.8 via_1600x480 ;
      VIA 344.9 35.36 via3_1600x480 ;
      VIA 344.9 35.36 via2_1600x480 ;
      VIA 344.9 35.36 via_1600x480 ;
      VIA 324.7 35.36 via3_1600x480 ;
      VIA 324.7 35.36 via2_1600x480 ;
      VIA 324.7 35.36 via_1600x480 ;
      VIA 304.5 35.36 via3_1600x480 ;
      VIA 304.5 35.36 via2_1600x480 ;
      VIA 304.5 35.36 via_1600x480 ;
      VIA 284.3 35.36 via3_1600x480 ;
      VIA 284.3 35.36 via2_1600x480 ;
      VIA 284.3 35.36 via_1600x480 ;
      VIA 264.1 35.36 via3_1600x480 ;
      VIA 264.1 35.36 via2_1600x480 ;
      VIA 264.1 35.36 via_1600x480 ;
      VIA 243.9 35.36 via3_1600x480 ;
      VIA 243.9 35.36 via2_1600x480 ;
      VIA 243.9 35.36 via_1600x480 ;
      VIA 223.7 35.36 via3_1600x480 ;
      VIA 223.7 35.36 via2_1600x480 ;
      VIA 223.7 35.36 via_1600x480 ;
      VIA 203.5 35.36 via3_1600x480 ;
      VIA 203.5 35.36 via2_1600x480 ;
      VIA 203.5 35.36 via_1600x480 ;
      VIA 183.3 35.36 via3_1600x480 ;
      VIA 183.3 35.36 via2_1600x480 ;
      VIA 183.3 35.36 via_1600x480 ;
      VIA 163.1 35.36 via3_1600x480 ;
      VIA 163.1 35.36 via2_1600x480 ;
      VIA 163.1 35.36 via_1600x480 ;
      VIA 142.9 35.36 via3_1600x480 ;
      VIA 142.9 35.36 via2_1600x480 ;
      VIA 142.9 35.36 via_1600x480 ;
      VIA 122.7 35.36 via3_1600x480 ;
      VIA 122.7 35.36 via2_1600x480 ;
      VIA 122.7 35.36 via_1600x480 ;
      VIA 102.5 35.36 via3_1600x480 ;
      VIA 102.5 35.36 via2_1600x480 ;
      VIA 102.5 35.36 via_1600x480 ;
      VIA 82.3 35.36 via3_1600x480 ;
      VIA 82.3 35.36 via2_1600x480 ;
      VIA 82.3 35.36 via_1600x480 ;
      VIA 62.1 35.36 via3_1600x480 ;
      VIA 62.1 35.36 via2_1600x480 ;
      VIA 62.1 35.36 via_1600x480 ;
      VIA 41.9 35.36 via3_1600x480 ;
      VIA 41.9 35.36 via2_1600x480 ;
      VIA 41.9 35.36 via_1600x480 ;
      VIA 21.7 35.36 via3_1600x480 ;
      VIA 21.7 35.36 via2_1600x480 ;
      VIA 21.7 35.36 via_1600x480 ;
      VIA 344.9 29.92 via3_1600x480 ;
      VIA 344.9 29.92 via2_1600x480 ;
      VIA 344.9 29.92 via_1600x480 ;
      VIA 324.7 29.92 via3_1600x480 ;
      VIA 324.7 29.92 via2_1600x480 ;
      VIA 324.7 29.92 via_1600x480 ;
      VIA 304.5 29.92 via3_1600x480 ;
      VIA 304.5 29.92 via2_1600x480 ;
      VIA 304.5 29.92 via_1600x480 ;
      VIA 284.3 29.92 via3_1600x480 ;
      VIA 284.3 29.92 via2_1600x480 ;
      VIA 284.3 29.92 via_1600x480 ;
      VIA 264.1 29.92 via3_1600x480 ;
      VIA 264.1 29.92 via2_1600x480 ;
      VIA 264.1 29.92 via_1600x480 ;
      VIA 243.9 29.92 via3_1600x480 ;
      VIA 243.9 29.92 via2_1600x480 ;
      VIA 243.9 29.92 via_1600x480 ;
      VIA 223.7 29.92 via3_1600x480 ;
      VIA 223.7 29.92 via2_1600x480 ;
      VIA 223.7 29.92 via_1600x480 ;
      VIA 203.5 29.92 via3_1600x480 ;
      VIA 203.5 29.92 via2_1600x480 ;
      VIA 203.5 29.92 via_1600x480 ;
      VIA 183.3 29.92 via3_1600x480 ;
      VIA 183.3 29.92 via2_1600x480 ;
      VIA 183.3 29.92 via_1600x480 ;
      VIA 163.1 29.92 via3_1600x480 ;
      VIA 163.1 29.92 via2_1600x480 ;
      VIA 163.1 29.92 via_1600x480 ;
      VIA 142.9 29.92 via3_1600x480 ;
      VIA 142.9 29.92 via2_1600x480 ;
      VIA 142.9 29.92 via_1600x480 ;
      VIA 122.7 29.92 via3_1600x480 ;
      VIA 122.7 29.92 via2_1600x480 ;
      VIA 122.7 29.92 via_1600x480 ;
      VIA 102.5 29.92 via3_1600x480 ;
      VIA 102.5 29.92 via2_1600x480 ;
      VIA 102.5 29.92 via_1600x480 ;
      VIA 82.3 29.92 via3_1600x480 ;
      VIA 82.3 29.92 via2_1600x480 ;
      VIA 82.3 29.92 via_1600x480 ;
      VIA 62.1 29.92 via3_1600x480 ;
      VIA 62.1 29.92 via2_1600x480 ;
      VIA 62.1 29.92 via_1600x480 ;
      VIA 41.9 29.92 via3_1600x480 ;
      VIA 41.9 29.92 via2_1600x480 ;
      VIA 41.9 29.92 via_1600x480 ;
      VIA 21.7 29.92 via3_1600x480 ;
      VIA 21.7 29.92 via2_1600x480 ;
      VIA 21.7 29.92 via_1600x480 ;
      VIA 344.9 24.48 via3_1600x480 ;
      VIA 344.9 24.48 via2_1600x480 ;
      VIA 344.9 24.48 via_1600x480 ;
      VIA 324.7 24.48 via3_1600x480 ;
      VIA 324.7 24.48 via2_1600x480 ;
      VIA 324.7 24.48 via_1600x480 ;
      VIA 304.5 24.48 via3_1600x480 ;
      VIA 304.5 24.48 via2_1600x480 ;
      VIA 304.5 24.48 via_1600x480 ;
      VIA 284.3 24.48 via3_1600x480 ;
      VIA 284.3 24.48 via2_1600x480 ;
      VIA 284.3 24.48 via_1600x480 ;
      VIA 264.1 24.48 via3_1600x480 ;
      VIA 264.1 24.48 via2_1600x480 ;
      VIA 264.1 24.48 via_1600x480 ;
      VIA 243.9 24.48 via3_1600x480 ;
      VIA 243.9 24.48 via2_1600x480 ;
      VIA 243.9 24.48 via_1600x480 ;
      VIA 223.7 24.48 via3_1600x480 ;
      VIA 223.7 24.48 via2_1600x480 ;
      VIA 223.7 24.48 via_1600x480 ;
      VIA 203.5 24.48 via3_1600x480 ;
      VIA 203.5 24.48 via2_1600x480 ;
      VIA 203.5 24.48 via_1600x480 ;
      VIA 183.3 24.48 via3_1600x480 ;
      VIA 183.3 24.48 via2_1600x480 ;
      VIA 183.3 24.48 via_1600x480 ;
      VIA 163.1 24.48 via3_1600x480 ;
      VIA 163.1 24.48 via2_1600x480 ;
      VIA 163.1 24.48 via_1600x480 ;
      VIA 142.9 24.48 via3_1600x480 ;
      VIA 142.9 24.48 via2_1600x480 ;
      VIA 142.9 24.48 via_1600x480 ;
      VIA 122.7 24.48 via3_1600x480 ;
      VIA 122.7 24.48 via2_1600x480 ;
      VIA 122.7 24.48 via_1600x480 ;
      VIA 102.5 24.48 via3_1600x480 ;
      VIA 102.5 24.48 via2_1600x480 ;
      VIA 102.5 24.48 via_1600x480 ;
      VIA 82.3 24.48 via3_1600x480 ;
      VIA 82.3 24.48 via2_1600x480 ;
      VIA 82.3 24.48 via_1600x480 ;
      VIA 62.1 24.48 via3_1600x480 ;
      VIA 62.1 24.48 via2_1600x480 ;
      VIA 62.1 24.48 via_1600x480 ;
      VIA 41.9 24.48 via3_1600x480 ;
      VIA 41.9 24.48 via2_1600x480 ;
      VIA 41.9 24.48 via_1600x480 ;
      VIA 21.7 24.48 via3_1600x480 ;
      VIA 21.7 24.48 via2_1600x480 ;
      VIA 21.7 24.48 via_1600x480 ;
      VIA 344.9 19.04 via3_1600x480 ;
      VIA 344.9 19.04 via2_1600x480 ;
      VIA 344.9 19.04 via_1600x480 ;
      VIA 324.7 19.04 via3_1600x480 ;
      VIA 324.7 19.04 via2_1600x480 ;
      VIA 324.7 19.04 via_1600x480 ;
      VIA 304.5 19.04 via3_1600x480 ;
      VIA 304.5 19.04 via2_1600x480 ;
      VIA 304.5 19.04 via_1600x480 ;
      VIA 284.3 19.04 via3_1600x480 ;
      VIA 284.3 19.04 via2_1600x480 ;
      VIA 284.3 19.04 via_1600x480 ;
      VIA 264.1 19.04 via3_1600x480 ;
      VIA 264.1 19.04 via2_1600x480 ;
      VIA 264.1 19.04 via_1600x480 ;
      VIA 243.9 19.04 via3_1600x480 ;
      VIA 243.9 19.04 via2_1600x480 ;
      VIA 243.9 19.04 via_1600x480 ;
      VIA 223.7 19.04 via3_1600x480 ;
      VIA 223.7 19.04 via2_1600x480 ;
      VIA 223.7 19.04 via_1600x480 ;
      VIA 203.5 19.04 via3_1600x480 ;
      VIA 203.5 19.04 via2_1600x480 ;
      VIA 203.5 19.04 via_1600x480 ;
      VIA 183.3 19.04 via3_1600x480 ;
      VIA 183.3 19.04 via2_1600x480 ;
      VIA 183.3 19.04 via_1600x480 ;
      VIA 163.1 19.04 via3_1600x480 ;
      VIA 163.1 19.04 via2_1600x480 ;
      VIA 163.1 19.04 via_1600x480 ;
      VIA 142.9 19.04 via3_1600x480 ;
      VIA 142.9 19.04 via2_1600x480 ;
      VIA 142.9 19.04 via_1600x480 ;
      VIA 122.7 19.04 via3_1600x480 ;
      VIA 122.7 19.04 via2_1600x480 ;
      VIA 122.7 19.04 via_1600x480 ;
      VIA 102.5 19.04 via3_1600x480 ;
      VIA 102.5 19.04 via2_1600x480 ;
      VIA 102.5 19.04 via_1600x480 ;
      VIA 82.3 19.04 via3_1600x480 ;
      VIA 82.3 19.04 via2_1600x480 ;
      VIA 82.3 19.04 via_1600x480 ;
      VIA 62.1 19.04 via3_1600x480 ;
      VIA 62.1 19.04 via2_1600x480 ;
      VIA 62.1 19.04 via_1600x480 ;
      VIA 41.9 19.04 via3_1600x480 ;
      VIA 41.9 19.04 via2_1600x480 ;
      VIA 41.9 19.04 via_1600x480 ;
      VIA 21.7 19.04 via3_1600x480 ;
      VIA 21.7 19.04 via2_1600x480 ;
      VIA 21.7 19.04 via_1600x480 ;
      VIA 344.9 13.6 via3_1600x480 ;
      VIA 344.9 13.6 via2_1600x480 ;
      VIA 344.9 13.6 via_1600x480 ;
      VIA 324.7 13.6 via3_1600x480 ;
      VIA 324.7 13.6 via2_1600x480 ;
      VIA 324.7 13.6 via_1600x480 ;
      VIA 304.5 13.6 via3_1600x480 ;
      VIA 304.5 13.6 via2_1600x480 ;
      VIA 304.5 13.6 via_1600x480 ;
      VIA 284.3 13.6 via3_1600x480 ;
      VIA 284.3 13.6 via2_1600x480 ;
      VIA 284.3 13.6 via_1600x480 ;
      VIA 264.1 13.6 via3_1600x480 ;
      VIA 264.1 13.6 via2_1600x480 ;
      VIA 264.1 13.6 via_1600x480 ;
      VIA 243.9 13.6 via3_1600x480 ;
      VIA 243.9 13.6 via2_1600x480 ;
      VIA 243.9 13.6 via_1600x480 ;
      VIA 223.7 13.6 via3_1600x480 ;
      VIA 223.7 13.6 via2_1600x480 ;
      VIA 223.7 13.6 via_1600x480 ;
      VIA 203.5 13.6 via3_1600x480 ;
      VIA 203.5 13.6 via2_1600x480 ;
      VIA 203.5 13.6 via_1600x480 ;
      VIA 183.3 13.6 via3_1600x480 ;
      VIA 183.3 13.6 via2_1600x480 ;
      VIA 183.3 13.6 via_1600x480 ;
      VIA 163.1 13.6 via3_1600x480 ;
      VIA 163.1 13.6 via2_1600x480 ;
      VIA 163.1 13.6 via_1600x480 ;
      VIA 142.9 13.6 via3_1600x480 ;
      VIA 142.9 13.6 via2_1600x480 ;
      VIA 142.9 13.6 via_1600x480 ;
      VIA 122.7 13.6 via3_1600x480 ;
      VIA 122.7 13.6 via2_1600x480 ;
      VIA 122.7 13.6 via_1600x480 ;
      VIA 102.5 13.6 via3_1600x480 ;
      VIA 102.5 13.6 via2_1600x480 ;
      VIA 102.5 13.6 via_1600x480 ;
      VIA 82.3 13.6 via3_1600x480 ;
      VIA 82.3 13.6 via2_1600x480 ;
      VIA 82.3 13.6 via_1600x480 ;
      VIA 62.1 13.6 via3_1600x480 ;
      VIA 62.1 13.6 via2_1600x480 ;
      VIA 62.1 13.6 via_1600x480 ;
      VIA 41.9 13.6 via3_1600x480 ;
      VIA 41.9 13.6 via2_1600x480 ;
      VIA 41.9 13.6 via_1600x480 ;
      VIA 21.7 13.6 via3_1600x480 ;
      VIA 21.7 13.6 via2_1600x480 ;
      VIA 21.7 13.6 via_1600x480 ;
      VIA 344.9 8.16 via3_1600x480 ;
      VIA 344.9 8.16 via2_1600x480 ;
      VIA 344.9 8.16 via_1600x480 ;
      VIA 324.7 8.16 via3_1600x480 ;
      VIA 324.7 8.16 via2_1600x480 ;
      VIA 324.7 8.16 via_1600x480 ;
      VIA 304.5 8.16 via3_1600x480 ;
      VIA 304.5 8.16 via2_1600x480 ;
      VIA 304.5 8.16 via_1600x480 ;
      VIA 284.3 8.16 via3_1600x480 ;
      VIA 284.3 8.16 via2_1600x480 ;
      VIA 284.3 8.16 via_1600x480 ;
      VIA 264.1 8.16 via3_1600x480 ;
      VIA 264.1 8.16 via2_1600x480 ;
      VIA 264.1 8.16 via_1600x480 ;
      VIA 243.9 8.16 via3_1600x480 ;
      VIA 243.9 8.16 via2_1600x480 ;
      VIA 243.9 8.16 via_1600x480 ;
      VIA 223.7 8.16 via3_1600x480 ;
      VIA 223.7 8.16 via2_1600x480 ;
      VIA 223.7 8.16 via_1600x480 ;
      VIA 203.5 8.16 via3_1600x480 ;
      VIA 203.5 8.16 via2_1600x480 ;
      VIA 203.5 8.16 via_1600x480 ;
      VIA 183.3 8.16 via3_1600x480 ;
      VIA 183.3 8.16 via2_1600x480 ;
      VIA 183.3 8.16 via_1600x480 ;
      VIA 163.1 8.16 via3_1600x480 ;
      VIA 163.1 8.16 via2_1600x480 ;
      VIA 163.1 8.16 via_1600x480 ;
      VIA 142.9 8.16 via3_1600x480 ;
      VIA 142.9 8.16 via2_1600x480 ;
      VIA 142.9 8.16 via_1600x480 ;
      VIA 122.7 8.16 via3_1600x480 ;
      VIA 122.7 8.16 via2_1600x480 ;
      VIA 122.7 8.16 via_1600x480 ;
      VIA 102.5 8.16 via3_1600x480 ;
      VIA 102.5 8.16 via2_1600x480 ;
      VIA 102.5 8.16 via_1600x480 ;
      VIA 82.3 8.16 via3_1600x480 ;
      VIA 82.3 8.16 via2_1600x480 ;
      VIA 82.3 8.16 via_1600x480 ;
      VIA 62.1 8.16 via3_1600x480 ;
      VIA 62.1 8.16 via2_1600x480 ;
      VIA 62.1 8.16 via_1600x480 ;
      VIA 41.9 8.16 via3_1600x480 ;
      VIA 41.9 8.16 via2_1600x480 ;
      VIA 41.9 8.16 via_1600x480 ;
      VIA 21.7 8.16 via3_1600x480 ;
      VIA 21.7 8.16 via2_1600x480 ;
      VIA 21.7 8.16 via_1600x480 ;
      VIA 344.9 2.72 via3_1600x480 ;
      VIA 344.9 2.72 via2_1600x480 ;
      VIA 344.9 2.72 via_1600x480 ;
      VIA 324.7 2.72 via3_1600x480 ;
      VIA 324.7 2.72 via2_1600x480 ;
      VIA 324.7 2.72 via_1600x480 ;
      VIA 304.5 2.72 via3_1600x480 ;
      VIA 304.5 2.72 via2_1600x480 ;
      VIA 304.5 2.72 via_1600x480 ;
      VIA 284.3 2.72 via3_1600x480 ;
      VIA 284.3 2.72 via2_1600x480 ;
      VIA 284.3 2.72 via_1600x480 ;
      VIA 264.1 2.72 via3_1600x480 ;
      VIA 264.1 2.72 via2_1600x480 ;
      VIA 264.1 2.72 via_1600x480 ;
      VIA 243.9 2.72 via3_1600x480 ;
      VIA 243.9 2.72 via2_1600x480 ;
      VIA 243.9 2.72 via_1600x480 ;
      VIA 223.7 2.72 via3_1600x480 ;
      VIA 223.7 2.72 via2_1600x480 ;
      VIA 223.7 2.72 via_1600x480 ;
      VIA 203.5 2.72 via3_1600x480 ;
      VIA 203.5 2.72 via2_1600x480 ;
      VIA 203.5 2.72 via_1600x480 ;
      VIA 183.3 2.72 via3_1600x480 ;
      VIA 183.3 2.72 via2_1600x480 ;
      VIA 183.3 2.72 via_1600x480 ;
      VIA 163.1 2.72 via3_1600x480 ;
      VIA 163.1 2.72 via2_1600x480 ;
      VIA 163.1 2.72 via_1600x480 ;
      VIA 142.9 2.72 via3_1600x480 ;
      VIA 142.9 2.72 via2_1600x480 ;
      VIA 142.9 2.72 via_1600x480 ;
      VIA 122.7 2.72 via3_1600x480 ;
      VIA 122.7 2.72 via2_1600x480 ;
      VIA 122.7 2.72 via_1600x480 ;
      VIA 102.5 2.72 via3_1600x480 ;
      VIA 102.5 2.72 via2_1600x480 ;
      VIA 102.5 2.72 via_1600x480 ;
      VIA 82.3 2.72 via3_1600x480 ;
      VIA 82.3 2.72 via2_1600x480 ;
      VIA 82.3 2.72 via_1600x480 ;
      VIA 62.1 2.72 via3_1600x480 ;
      VIA 62.1 2.72 via2_1600x480 ;
      VIA 62.1 2.72 via_1600x480 ;
      VIA 41.9 2.72 via3_1600x480 ;
      VIA 41.9 2.72 via2_1600x480 ;
      VIA 41.9 2.72 via_1600x480 ;
      VIA 21.7 2.72 via3_1600x480 ;
      VIA 21.7 2.72 via2_1600x480 ;
      VIA 21.7 2.72 via_1600x480 ;
      LAYER met5 ;
        RECT  0 184.98 349.6 186.58 ;
        RECT  0 164.78 349.6 166.38 ;
        RECT  0 144.58 349.6 146.18 ;
        RECT  0 124.38 349.6 125.98 ;
        RECT  0 104.18 349.6 105.78 ;
        RECT  0 83.98 349.6 85.58 ;
        RECT  0 63.78 349.6 65.38 ;
        RECT  0 43.58 349.6 45.18 ;
        RECT  0 23.38 349.6 24.98 ;
      LAYER met4 ;
        RECT  344.1 2.48 345.7 198.8 ;
        RECT  323.9 2.48 325.5 198.8 ;
        RECT  303.7 2.48 305.3 198.8 ;
        RECT  283.5 2.48 285.1 198.8 ;
        RECT  263.3 2.48 264.9 198.8 ;
        RECT  243.1 2.48 244.7 198.8 ;
        RECT  222.9 2.48 224.5 198.8 ;
        RECT  202.7 2.48 204.3 198.8 ;
        RECT  182.5 2.48 184.1 198.8 ;
        RECT  162.3 2.48 163.9 198.8 ;
        RECT  142.1 2.48 143.7 198.8 ;
        RECT  121.9 2.48 123.5 198.8 ;
        RECT  101.7 2.48 103.3 198.8 ;
        RECT  81.5 2.48 83.1 198.8 ;
        RECT  61.3 2.48 62.9 198.8 ;
        RECT  41.1 2.48 42.7 198.8 ;
        RECT  20.9 2.48 22.5 198.8 ;
      LAYER met1 ;
        RECT  0 198.32 349.6 198.8 ;
        RECT  0 192.88 349.6 193.36 ;
        RECT  0 187.44 349.6 187.92 ;
        RECT  0 182 349.6 182.48 ;
        RECT  0 176.56 349.6 177.04 ;
        RECT  0 171.12 349.6 171.6 ;
        RECT  0 165.68 349.6 166.16 ;
        RECT  0 160.24 349.6 160.72 ;
        RECT  0 154.8 349.6 155.28 ;
        RECT  0 149.36 349.6 149.84 ;
        RECT  0 143.92 349.6 144.4 ;
        RECT  0 138.48 349.6 138.96 ;
        RECT  0 133.04 349.6 133.52 ;
        RECT  0 127.6 349.6 128.08 ;
        RECT  0 122.16 349.6 122.64 ;
        RECT  0 116.72 349.6 117.2 ;
        RECT  0 111.28 349.6 111.76 ;
        RECT  0 105.84 349.6 106.32 ;
        RECT  0 100.4 349.6 100.88 ;
        RECT  0 94.96 349.6 95.44 ;
        RECT  0 89.52 349.6 90 ;
        RECT  0 84.08 349.6 84.56 ;
        RECT  0 78.64 349.6 79.12 ;
        RECT  0 73.2 349.6 73.68 ;
        RECT  0 67.76 349.6 68.24 ;
        RECT  0 62.32 349.6 62.8 ;
        RECT  0 56.88 349.6 57.36 ;
        RECT  0 51.44 349.6 51.92 ;
        RECT  0 46 349.6 46.48 ;
        RECT  0 40.56 349.6 41.04 ;
        RECT  0 35.12 349.6 35.6 ;
        RECT  0 29.68 349.6 30.16 ;
        RECT  0 24.24 349.6 24.72 ;
        RECT  0 18.8 349.6 19.28 ;
        RECT  0 13.36 349.6 13.84 ;
        RECT  0 7.92 349.6 8.4 ;
        RECT  0 2.48 349.6 2.96 ;
    END
  END VSS
  PIN bl_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 61.39 0.8 61.69 ;
    END
  END bl_address[0]
  PIN bl_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  321.24 201.515 321.38 202 ;
    END
  END bl_address[1]
  PIN bl_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  71 201.515 71.14 202 ;
    END
  END bl_address[2]
  PIN bl_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  249.48 0 249.62 0.485 ;
    END
  END bl_address[3]
  PIN bl_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  153.8 201.515 153.94 202 ;
    END
  END bl_address[4]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  270.64 0 270.78 0.485 ;
    END
  END clk
  PIN data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  145.52 0 145.66 0.485 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 91.31 0.8 91.61 ;
    END
  END enable
  PIN gfpga_pad_GPIO_PAD[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  133.56 201.515 133.7 202 ;
    END
  END gfpga_pad_GPIO_PAD[0]
  PIN gfpga_pad_GPIO_PAD[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  229.24 0 229.38 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[10]
  PIN gfpga_pad_GPIO_PAD[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  290.88 0 291.02 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[11]
  PIN gfpga_pad_GPIO_PAD[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  351.2 156.59 352 156.89 ;
    END
  END gfpga_pad_GPIO_PAD[12]
  PIN gfpga_pad_GPIO_PAD[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  49.84 201.515 49.98 202 ;
    END
  END gfpga_pad_GPIO_PAD[13]
  PIN gfpga_pad_GPIO_PAD[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 122.59 0.8 122.89 ;
    END
  END gfpga_pad_GPIO_PAD[14]
  PIN gfpga_pad_GPIO_PAD[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  351.2 125.31 352 125.61 ;
    END
  END gfpga_pad_GPIO_PAD[15]
  PIN gfpga_pad_GPIO_PAD[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  186.92 0 187.06 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[16]
  PIN gfpga_pad_GPIO_PAD[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  278.92 201.515 279.06 202 ;
    END
  END gfpga_pad_GPIO_PAD[17]
  PIN gfpga_pad_GPIO_PAD[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 201.515 29.74 202 ;
    END
  END gfpga_pad_GPIO_PAD[18]
  PIN gfpga_pad_GPIO_PAD[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  112.4 201.515 112.54 202 ;
    END
  END gfpga_pad_GPIO_PAD[19]
  PIN gfpga_pad_GPIO_PAD[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  300.08 201.515 300.22 202 ;
    END
  END gfpga_pad_GPIO_PAD[1]
  PIN gfpga_pad_GPIO_PAD[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  237.52 201.515 237.66 202 ;
    END
  END gfpga_pad_GPIO_PAD[20]
  PIN gfpga_pad_GPIO_PAD[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 183.79 0.8 184.09 ;
    END
  END gfpga_pad_GPIO_PAD[21]
  PIN gfpga_pad_GPIO_PAD[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  351.2 64.11 352 64.41 ;
    END
  END gfpga_pad_GPIO_PAD[22]
  PIN gfpga_pad_GPIO_PAD[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 30.11 0.8 30.41 ;
    END
  END gfpga_pad_GPIO_PAD[23]
  PIN gfpga_pad_GPIO_PAD[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  8.44 201.515 8.58 202 ;
    END
  END gfpga_pad_GPIO_PAD[24]
  PIN gfpga_pad_GPIO_PAD[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 0 20.54 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[25]
  PIN gfpga_pad_GPIO_PAD[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  0.16 0 0.3 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[26]
  PIN gfpga_pad_GPIO_PAD[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  216.36 201.515 216.5 202 ;
    END
  END gfpga_pad_GPIO_PAD[27]
  PIN gfpga_pad_GPIO_PAD[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  351.2 94.03 352 94.33 ;
    END
  END gfpga_pad_GPIO_PAD[28]
  PIN gfpga_pad_GPIO_PAD[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  82.96 0 83.1 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[29]
  PIN gfpga_pad_GPIO_PAD[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  351.2 32.83 352 33.13 ;
    END
  END gfpga_pad_GPIO_PAD[2]
  PIN gfpga_pad_GPIO_PAD[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  208.08 0 208.22 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[30]
  PIN gfpga_pad_GPIO_PAD[31]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  258.68 201.515 258.82 202 ;
    END
  END gfpga_pad_GPIO_PAD[31]
  PIN gfpga_pad_GPIO_PAD[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  312.04 0 312.18 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[3]
  PIN gfpga_pad_GPIO_PAD[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  41.56 0 41.7 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[4]
  PIN gfpga_pad_GPIO_PAD[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  61.8 0 61.94 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[5]
  PIN gfpga_pad_GPIO_PAD[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  104.12 0 104.26 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[6]
  PIN gfpga_pad_GPIO_PAD[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  333.2 0 333.34 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[7]
  PIN gfpga_pad_GPIO_PAD[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  124.36 0 124.5 0.485 ;
    END
  END gfpga_pad_GPIO_PAD[8]
  PIN gfpga_pad_GPIO_PAD[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  351.2 186.51 352 186.81 ;
    END
  END gfpga_pad_GPIO_PAD[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  341.48 201.515 341.62 202 ;
    END
  END reset
  PIN set
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.96 201.515 175.1 202 ;
    END
  END set
  PIN wl_address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  196.12 201.515 196.26 202 ;
    END
  END wl_address[0]
  PIN wl_address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  166.68 0 166.82 0.485 ;
    END
  END wl_address[1]
  PIN wl_address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 153.87 0.8 154.17 ;
    END
  END wl_address[2]
  PIN wl_address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.16 201.515 92.3 202 ;
    END
  END wl_address[3]
  PIN wl_address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  351.2 1.55 352 1.85 ;
    END
  END wl_address[4]
  OBS
    LAYER li1 ;
    RECT  0 0 352.05 202 ;
    LAYER met1 ;
    RECT  0 0 352.05 202 ;
    LAYER via ;
    RECT  0 0 352.05 202 ;
    LAYER met2 ;
    RECT  0 0 352.05 202 ;
    LAYER via2 ;
    RECT  0 0 352.05 202 ;
    LAYER met3 ;
    RECT  0 0 352.05 202 ;
    LAYER via3 ;
    RECT  0 0 352.05 202 ;
    LAYER met4 ;
    RECT  0 0 352.05 202 ;
    LAYER via4 ;
    RECT  0 0 352.05 202 ;
    LAYER met5 ;
    RECT  0 0 352.05 202 ;
  END
END test_lut_inst
END LIBRARY
