VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wl_driver
  CLASS BLOCK ;
  FOREIGN wl_driver ;
  ORIGIN 12.500 4.430 ;
  SIZE 124.110 BY 8.645 ;
  PIN OUT[31]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 110.900 -2.015 111.155 0.345 ;
        RECT 110.955 -2.685 111.155 -2.015 ;
        RECT 110.900 -3.565 111.155 -2.685 ;
    END
  END OUT[31]
  PIN OUT[30]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 107.540 -2.015 107.795 0.345 ;
        RECT 107.595 -2.685 107.795 -2.015 ;
        RECT 107.540 -3.565 107.795 -2.685 ;
    END
  END OUT[30]
  PIN OUT[29]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 104.180 -2.015 104.435 0.345 ;
        RECT 104.235 -2.685 104.435 -2.015 ;
        RECT 104.180 -3.565 104.435 -2.685 ;
    END
  END OUT[29]
  PIN OUT[28]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 100.820 -2.015 101.075 0.345 ;
        RECT 100.875 -2.685 101.075 -2.015 ;
        RECT 100.820 -3.565 101.075 -2.685 ;
    END
  END OUT[28]
  PIN OUT[27]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 97.460 -2.015 97.715 0.345 ;
        RECT 97.515 -2.685 97.715 -2.015 ;
        RECT 97.460 -3.565 97.715 -2.685 ;
    END
  END OUT[27]
  PIN OUT[26]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 94.100 -2.015 94.355 0.345 ;
        RECT 94.155 -2.685 94.355 -2.015 ;
        RECT 94.100 -3.565 94.355 -2.685 ;
    END
  END OUT[26]
  PIN OUT[25]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 90.740 -2.015 90.995 0.345 ;
        RECT 90.795 -2.685 90.995 -2.015 ;
        RECT 90.740 -3.565 90.995 -2.685 ;
    END
  END OUT[25]
  PIN OUT[24]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 87.380 -2.015 87.635 0.345 ;
        RECT 87.435 -2.685 87.635 -2.015 ;
        RECT 87.380 -3.565 87.635 -2.685 ;
    END
  END OUT[24]
  PIN OUT[23]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 84.020 -2.015 84.275 0.345 ;
        RECT 84.075 -2.685 84.275 -2.015 ;
        RECT 84.020 -3.565 84.275 -2.685 ;
    END
  END OUT[23]
  PIN OUT[22]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 80.660 -2.015 80.915 0.345 ;
        RECT 80.715 -2.685 80.915 -2.015 ;
        RECT 80.660 -3.565 80.915 -2.685 ;
    END
  END OUT[22]
  PIN OUT[21]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 77.300 -2.015 77.555 0.345 ;
        RECT 77.355 -2.685 77.555 -2.015 ;
        RECT 77.300 -3.565 77.555 -2.685 ;
    END
  END OUT[21]
  PIN OUT[20]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 73.940 -2.015 74.195 0.345 ;
        RECT 73.995 -2.685 74.195 -2.015 ;
        RECT 73.940 -3.565 74.195 -2.685 ;
    END
  END OUT[20]
  PIN OUT[19]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 70.580 -2.015 70.835 0.345 ;
        RECT 70.635 -2.685 70.835 -2.015 ;
        RECT 70.580 -3.565 70.835 -2.685 ;
    END
  END OUT[19]
  PIN OUT[18]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 67.220 -2.015 67.475 0.345 ;
        RECT 67.275 -2.685 67.475 -2.015 ;
        RECT 67.220 -3.565 67.475 -2.685 ;
    END
  END OUT[18]
  PIN OUT[17]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 63.860 -2.015 64.115 0.345 ;
        RECT 63.915 -2.685 64.115 -2.015 ;
        RECT 63.860 -3.565 64.115 -2.685 ;
    END
  END OUT[17]
  PIN OUT[16]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 60.500 -2.015 60.755 0.345 ;
        RECT 60.555 -2.685 60.755 -2.015 ;
        RECT 60.500 -3.565 60.755 -2.685 ;
    END
  END OUT[16]
  PIN OUT[15]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 57.140 -2.015 57.395 0.345 ;
        RECT 57.195 -2.685 57.395 -2.015 ;
        RECT 57.140 -3.565 57.395 -2.685 ;
    END
  END OUT[15]
  PIN OUT[14]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 53.780 -2.015 54.035 0.345 ;
        RECT 53.835 -2.685 54.035 -2.015 ;
        RECT 53.780 -3.565 54.035 -2.685 ;
    END
  END OUT[14]
  PIN OUT[13]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 50.420 -2.015 50.675 0.345 ;
        RECT 50.475 -2.685 50.675 -2.015 ;
        RECT 50.420 -3.565 50.675 -2.685 ;
    END
  END OUT[13]
  PIN OUT[12]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 47.060 -2.015 47.315 0.345 ;
        RECT 47.115 -2.685 47.315 -2.015 ;
        RECT 47.060 -3.565 47.315 -2.685 ;
    END
  END OUT[12]
  PIN OUT[11]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 43.700 -2.015 43.955 0.345 ;
        RECT 43.755 -2.685 43.955 -2.015 ;
        RECT 43.700 -3.565 43.955 -2.685 ;
    END
  END OUT[11]
  PIN OUT[10]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 40.340 -2.015 40.595 0.345 ;
        RECT 40.395 -2.685 40.595 -2.015 ;
        RECT 40.340 -3.565 40.595 -2.685 ;
    END
  END OUT[10]
  PIN OUT[9]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 36.980 -2.015 37.235 0.345 ;
        RECT 37.035 -2.685 37.235 -2.015 ;
        RECT 36.980 -3.565 37.235 -2.685 ;
    END
  END OUT[9]
  PIN OUT[8]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 33.620 -2.015 33.875 0.345 ;
        RECT 33.675 -2.685 33.875 -2.015 ;
        RECT 33.620 -3.565 33.875 -2.685 ;
    END
  END OUT[8]
  PIN OUT[7]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 30.260 -2.015 30.515 0.345 ;
        RECT 30.315 -2.685 30.515 -2.015 ;
        RECT 30.260 -3.565 30.515 -2.685 ;
    END
  END OUT[7]
  PIN OUT[6]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 26.900 -2.015 27.155 0.345 ;
        RECT 26.955 -2.685 27.155 -2.015 ;
        RECT 26.900 -3.565 27.155 -2.685 ;
    END
  END OUT[6]
  PIN OUT[5]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 23.540 -2.015 23.795 0.345 ;
        RECT 23.595 -2.685 23.795 -2.015 ;
        RECT 23.540 -3.565 23.795 -2.685 ;
    END
  END OUT[5]
  PIN OUT[4]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 20.180 -2.015 20.435 0.345 ;
        RECT 20.235 -2.685 20.435 -2.015 ;
        RECT 20.180 -3.565 20.435 -2.685 ;
    END
  END OUT[4]
  PIN OUT[3]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 16.820 -2.015 17.075 0.345 ;
        RECT 16.875 -2.685 17.075 -2.015 ;
        RECT 16.820 -3.565 17.075 -2.685 ;
    END
  END OUT[3]
  PIN OUT[2]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 13.460 -2.015 13.715 0.345 ;
        RECT 13.515 -2.685 13.715 -2.015 ;
        RECT 13.460 -3.565 13.715 -2.685 ;
    END
  END OUT[2]
  PIN OUT[1]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 10.100 -2.015 10.355 0.345 ;
        RECT 10.155 -2.685 10.355 -2.015 ;
        RECT 10.100 -3.565 10.355 -2.685 ;
    END
  END OUT[1]
  PIN OUT[0]
    ANTENNADIFFAREA 0.641250 ;
    PORT
      LAYER li1 ;
        RECT 6.740 -2.015 6.995 0.345 ;
        RECT 6.795 -2.685 6.995 -2.015 ;
        RECT 6.740 -3.565 6.995 -2.685 ;
    END
  END OUT[0]
  PIN VRO
    ANTENNADIFFAREA 0.665800 ;
    PORT
      LAYER li1 ;
        RECT -2.620 1.290 -1.255 1.700 ;
        RECT -2.620 0.245 -0.590 1.290 ;
      LAYER mcon ;
        RECT -2.590 0.325 -2.420 0.495 ;
        RECT -2.230 0.325 -2.060 0.495 ;
        RECT -1.870 0.325 -1.700 0.495 ;
        RECT -1.510 0.325 -1.340 0.495 ;
        RECT -1.150 0.325 -0.980 0.495 ;
        RECT -0.790 0.325 -0.620 0.495 ;
      LAYER met1 ;
        RECT -3.360 0.550 0.000 0.555 ;
        RECT -12.500 0.190 0.000 0.550 ;
        RECT -3.360 0.185 0.000 0.190 ;
    END
  END VRO
  PIN VHV
    ANTENNADIFFAREA 0.978150 ;
    PORT
      LAYER nwell ;
        RECT -3.690 -2.255 0.330 2.115 ;
      LAYER li1 ;
        RECT -3.360 -0.155 -0.635 0.015 ;
        RECT -2.530 -1.430 -0.560 -0.385 ;
        RECT -2.530 -1.860 -1.085 -1.430 ;
      LAYER mcon ;
        RECT -3.205 -0.155 -3.035 0.015 ;
        RECT -2.725 -0.155 -2.555 0.015 ;
        RECT -2.245 -0.155 -2.075 0.015 ;
        RECT -1.765 -0.155 -1.595 0.015 ;
        RECT -1.285 -0.155 -1.115 0.015 ;
        RECT -0.805 -0.155 -0.635 0.015 ;
        RECT -2.530 -0.635 -2.360 -0.465 ;
        RECT -2.170 -0.635 -2.000 -0.465 ;
        RECT -1.810 -0.635 -1.640 -0.465 ;
        RECT -1.450 -0.635 -1.280 -0.465 ;
        RECT -1.090 -0.635 -0.920 -0.465 ;
        RECT -0.730 -0.635 -0.560 -0.465 ;
      LAYER met1 ;
        RECT -3.360 -0.170 -0.540 0.045 ;
        RECT -12.500 -0.325 -0.540 -0.170 ;
        RECT -12.500 -0.530 0.000 -0.325 ;
        RECT -3.360 -0.695 0.000 -0.530 ;
    END
  END VHV
  PIN MODE
    ANTENNAGATEAREA 2.295000 ;
    PORT
      LAYER li1 ;
        RECT -2.845 1.975 -1.565 2.175 ;
        RECT -2.725 1.880 -1.565 1.975 ;
        RECT -2.845 -2.635 -2.055 -2.390 ;
      LAYER mcon ;
        RECT -2.490 1.955 -2.320 2.125 ;
        RECT -2.490 -2.565 -2.320 -2.395 ;
      LAYER met1 ;
        RECT -2.660 1.760 -2.190 2.290 ;
        RECT -2.750 -2.770 -2.130 -2.240 ;
      LAYER via ;
        RECT -2.545 1.905 -2.265 2.185 ;
        RECT -2.545 -2.625 -2.265 -2.345 ;
      LAYER met2 ;
        RECT -2.660 -4.360 -2.190 2.290 ;
    END
  END MODE
  PIN G_ENABLE
    ANTENNAGATEAREA 2.250000 ;
    PORT
      LAYER li1 ;
        RECT -0.855 2.275 -0.580 2.840 ;
        RECT -1.085 1.460 -0.580 2.275 ;
        RECT -0.915 -2.185 -0.550 -1.600 ;
        RECT -1.085 -2.515 -0.495 -2.185 ;
        RECT -0.915 -2.980 -0.550 -2.515 ;
      LAYER mcon ;
        RECT -0.920 1.985 -0.750 2.155 ;
        RECT -0.860 -2.435 -0.690 -2.265 ;
      LAYER met1 ;
        RECT -1.040 1.810 1.060 2.310 ;
        RECT 0.620 -1.410 1.060 1.810 ;
        RECT -3.360 -1.650 1.060 -1.410 ;
        RECT -0.940 -2.600 -0.540 -1.650 ;
        RECT 0.620 -2.590 1.060 -1.650 ;
      LAYER via ;
        RECT 0.695 -2.495 0.975 -2.215 ;
      LAYER met2 ;
        RECT 0.620 -4.430 1.090 -2.100 ;
    END
  END G_ENABLE
  PIN DATA
    ANTENNAGATEAREA 36.000000 ;
    PORT
      LAYER li1 ;
        RECT 6.205 -2.185 6.570 -1.600 ;
        RECT 9.565 -2.185 9.930 -1.600 ;
        RECT 12.925 -2.185 13.290 -1.600 ;
        RECT 16.285 -2.185 16.650 -1.600 ;
        RECT 19.645 -2.185 20.010 -1.600 ;
        RECT 23.005 -2.185 23.370 -1.600 ;
        RECT 26.365 -2.185 26.730 -1.600 ;
        RECT 29.725 -2.185 30.090 -1.600 ;
        RECT 33.085 -2.185 33.450 -1.600 ;
        RECT 36.445 -2.185 36.810 -1.600 ;
        RECT 39.805 -2.185 40.170 -1.600 ;
        RECT 43.165 -2.185 43.530 -1.600 ;
        RECT 46.525 -2.185 46.890 -1.600 ;
        RECT 49.885 -2.185 50.250 -1.600 ;
        RECT 53.245 -2.185 53.610 -1.600 ;
        RECT 56.605 -2.185 56.970 -1.600 ;
        RECT 59.965 -2.185 60.330 -1.600 ;
        RECT 63.325 -2.185 63.690 -1.600 ;
        RECT 66.685 -2.185 67.050 -1.600 ;
        RECT 70.045 -2.185 70.410 -1.600 ;
        RECT 73.405 -2.185 73.770 -1.600 ;
        RECT 76.765 -2.185 77.130 -1.600 ;
        RECT 80.125 -2.185 80.490 -1.600 ;
        RECT 83.485 -2.185 83.850 -1.600 ;
        RECT 86.845 -2.185 87.210 -1.600 ;
        RECT 90.205 -2.185 90.570 -1.600 ;
        RECT 93.565 -2.185 93.930 -1.600 ;
        RECT 96.925 -2.185 97.290 -1.600 ;
        RECT 100.285 -2.185 100.650 -1.600 ;
        RECT 103.645 -2.185 104.010 -1.600 ;
        RECT 107.005 -2.185 107.370 -1.600 ;
        RECT 110.365 -2.185 110.730 -1.600 ;
        RECT 6.035 -2.515 6.625 -2.185 ;
        RECT 9.395 -2.515 9.985 -2.185 ;
        RECT 12.755 -2.515 13.345 -2.185 ;
        RECT 16.115 -2.515 16.705 -2.185 ;
        RECT 19.475 -2.515 20.065 -2.185 ;
        RECT 22.835 -2.515 23.425 -2.185 ;
        RECT 26.195 -2.515 26.785 -2.185 ;
        RECT 29.555 -2.515 30.145 -2.185 ;
        RECT 32.915 -2.515 33.505 -2.185 ;
        RECT 36.275 -2.515 36.865 -2.185 ;
        RECT 39.635 -2.515 40.225 -2.185 ;
        RECT 42.995 -2.515 43.585 -2.185 ;
        RECT 46.355 -2.515 46.945 -2.185 ;
        RECT 49.715 -2.515 50.305 -2.185 ;
        RECT 53.075 -2.515 53.665 -2.185 ;
        RECT 56.435 -2.515 57.025 -2.185 ;
        RECT 59.795 -2.515 60.385 -2.185 ;
        RECT 63.155 -2.515 63.745 -2.185 ;
        RECT 66.515 -2.515 67.105 -2.185 ;
        RECT 69.875 -2.515 70.465 -2.185 ;
        RECT 73.235 -2.515 73.825 -2.185 ;
        RECT 76.595 -2.515 77.185 -2.185 ;
        RECT 79.955 -2.515 80.545 -2.185 ;
        RECT 83.315 -2.515 83.905 -2.185 ;
        RECT 86.675 -2.515 87.265 -2.185 ;
        RECT 90.035 -2.515 90.625 -2.185 ;
        RECT 93.395 -2.515 93.985 -2.185 ;
        RECT 96.755 -2.515 97.345 -2.185 ;
        RECT 100.115 -2.515 100.705 -2.185 ;
        RECT 103.475 -2.515 104.065 -2.185 ;
        RECT 106.835 -2.515 107.425 -2.185 ;
        RECT 110.195 -2.515 110.785 -2.185 ;
        RECT 6.205 -2.980 6.570 -2.515 ;
        RECT 9.565 -2.980 9.930 -2.515 ;
        RECT 12.925 -2.980 13.290 -2.515 ;
        RECT 16.285 -2.980 16.650 -2.515 ;
        RECT 19.645 -2.980 20.010 -2.515 ;
        RECT 23.005 -2.980 23.370 -2.515 ;
        RECT 26.365 -2.980 26.730 -2.515 ;
        RECT 29.725 -2.980 30.090 -2.515 ;
        RECT 33.085 -2.980 33.450 -2.515 ;
        RECT 36.445 -2.980 36.810 -2.515 ;
        RECT 39.805 -2.980 40.170 -2.515 ;
        RECT 43.165 -2.980 43.530 -2.515 ;
        RECT 46.525 -2.980 46.890 -2.515 ;
        RECT 49.885 -2.980 50.250 -2.515 ;
        RECT 53.245 -2.980 53.610 -2.515 ;
        RECT 56.605 -2.980 56.970 -2.515 ;
        RECT 59.965 -2.980 60.330 -2.515 ;
        RECT 63.325 -2.980 63.690 -2.515 ;
        RECT 66.685 -2.980 67.050 -2.515 ;
        RECT 70.045 -2.980 70.410 -2.515 ;
        RECT 73.405 -2.980 73.770 -2.515 ;
        RECT 76.765 -2.980 77.130 -2.515 ;
        RECT 80.125 -2.980 80.490 -2.515 ;
        RECT 83.485 -2.980 83.850 -2.515 ;
        RECT 86.845 -2.980 87.210 -2.515 ;
        RECT 90.205 -2.980 90.570 -2.515 ;
        RECT 93.565 -2.980 93.930 -2.515 ;
        RECT 96.925 -2.980 97.290 -2.515 ;
        RECT 100.285 -2.980 100.650 -2.515 ;
        RECT 103.645 -2.980 104.010 -2.515 ;
        RECT 107.005 -2.980 107.370 -2.515 ;
        RECT 110.365 -2.980 110.730 -2.515 ;
      LAYER mcon ;
        RECT 6.260 -2.435 6.430 -2.265 ;
        RECT 9.620 -2.435 9.790 -2.265 ;
        RECT 12.980 -2.435 13.150 -2.265 ;
        RECT 16.340 -2.435 16.510 -2.265 ;
        RECT 19.700 -2.435 19.870 -2.265 ;
        RECT 23.060 -2.435 23.230 -2.265 ;
        RECT 26.420 -2.435 26.590 -2.265 ;
        RECT 29.780 -2.435 29.950 -2.265 ;
        RECT 33.140 -2.435 33.310 -2.265 ;
        RECT 36.500 -2.435 36.670 -2.265 ;
        RECT 39.860 -2.435 40.030 -2.265 ;
        RECT 43.220 -2.435 43.390 -2.265 ;
        RECT 46.580 -2.435 46.750 -2.265 ;
        RECT 49.940 -2.435 50.110 -2.265 ;
        RECT 53.300 -2.435 53.470 -2.265 ;
        RECT 56.660 -2.435 56.830 -2.265 ;
        RECT 60.020 -2.435 60.190 -2.265 ;
        RECT 63.380 -2.435 63.550 -2.265 ;
        RECT 66.740 -2.435 66.910 -2.265 ;
        RECT 70.100 -2.435 70.270 -2.265 ;
        RECT 73.460 -2.435 73.630 -2.265 ;
        RECT 76.820 -2.435 76.990 -2.265 ;
        RECT 80.180 -2.435 80.350 -2.265 ;
        RECT 83.540 -2.435 83.710 -2.265 ;
        RECT 86.900 -2.435 87.070 -2.265 ;
        RECT 90.260 -2.435 90.430 -2.265 ;
        RECT 93.620 -2.435 93.790 -2.265 ;
        RECT 96.980 -2.435 97.150 -2.265 ;
        RECT 100.340 -2.435 100.510 -2.265 ;
        RECT 103.700 -2.435 103.870 -2.265 ;
        RECT 107.060 -2.435 107.230 -2.265 ;
        RECT 110.420 -2.435 110.590 -2.265 ;
      LAYER met1 ;
        RECT 1.910 -1.650 111.280 -1.410 ;
        RECT 1.910 -2.840 2.530 -1.650 ;
        RECT 6.180 -2.600 6.580 -1.650 ;
        RECT 9.540 -2.600 9.940 -1.650 ;
        RECT 12.900 -2.600 13.300 -1.650 ;
        RECT 16.260 -2.600 16.660 -1.650 ;
        RECT 19.620 -2.600 20.020 -1.650 ;
        RECT 22.980 -2.600 23.380 -1.650 ;
        RECT 26.340 -2.600 26.740 -1.650 ;
        RECT 29.700 -2.600 30.100 -1.650 ;
        RECT 33.060 -2.600 33.460 -1.650 ;
        RECT 36.420 -2.600 36.820 -1.650 ;
        RECT 39.780 -2.600 40.180 -1.650 ;
        RECT 43.140 -2.600 43.540 -1.650 ;
        RECT 46.500 -2.600 46.900 -1.650 ;
        RECT 49.860 -2.600 50.260 -1.650 ;
        RECT 53.220 -2.600 53.620 -1.650 ;
        RECT 56.580 -2.600 56.980 -1.650 ;
        RECT 59.940 -2.600 60.340 -1.650 ;
        RECT 63.300 -2.600 63.700 -1.650 ;
        RECT 66.660 -2.600 67.060 -1.650 ;
        RECT 70.020 -2.600 70.420 -1.650 ;
        RECT 73.380 -2.600 73.780 -1.650 ;
        RECT 76.740 -2.600 77.140 -1.650 ;
        RECT 80.100 -2.600 80.500 -1.650 ;
        RECT 83.460 -2.600 83.860 -1.650 ;
        RECT 86.820 -2.600 87.220 -1.650 ;
        RECT 90.180 -2.600 90.580 -1.650 ;
        RECT 93.540 -2.600 93.940 -1.650 ;
        RECT 96.900 -2.600 97.300 -1.650 ;
        RECT 100.260 -2.600 100.660 -1.650 ;
        RECT 103.620 -2.600 104.020 -1.650 ;
        RECT 106.980 -2.600 107.380 -1.650 ;
        RECT 110.340 -2.600 110.740 -1.650 ;
      LAYER via ;
        RECT 2.085 -2.665 2.365 -2.385 ;
      LAYER met2 ;
        RECT 2.000 -4.430 2.470 -2.310 ;
    END
  END DATA
  PIN SEL[0]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 4.275 -2.635 5.065 -2.390 ;
      LAYER mcon ;
        RECT 4.630 -2.565 4.800 -2.395 ;
      LAYER met1 ;
        RECT 4.370 -2.770 4.990 -2.240 ;
      LAYER via ;
        RECT 4.575 -2.625 4.855 -2.345 ;
      LAYER met2 ;
        RECT 4.460 -4.360 4.930 -2.240 ;
    END
  END SEL[0]
  PIN SEL[1]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 7.635 -2.635 8.425 -2.390 ;
      LAYER mcon ;
        RECT 7.990 -2.565 8.160 -2.395 ;
      LAYER met1 ;
        RECT 7.730 -2.770 8.350 -2.240 ;
      LAYER via ;
        RECT 7.935 -2.625 8.215 -2.345 ;
      LAYER met2 ;
        RECT 7.820 -4.360 8.290 -2.240 ;
    END
  END SEL[1]
  PIN SEL[2]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 10.995 -2.635 11.785 -2.390 ;
      LAYER mcon ;
        RECT 11.350 -2.565 11.520 -2.395 ;
      LAYER met1 ;
        RECT 11.090 -2.770 11.710 -2.240 ;
      LAYER via ;
        RECT 11.295 -2.625 11.575 -2.345 ;
      LAYER met2 ;
        RECT 11.180 -4.360 11.650 -2.240 ;
    END
  END SEL[2]
  PIN SEL[3]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 14.355 -2.635 15.145 -2.390 ;
      LAYER mcon ;
        RECT 14.710 -2.565 14.880 -2.395 ;
      LAYER met1 ;
        RECT 14.450 -2.770 15.070 -2.240 ;
      LAYER via ;
        RECT 14.655 -2.625 14.935 -2.345 ;
      LAYER met2 ;
        RECT 14.540 -4.360 15.010 -2.240 ;
    END
  END SEL[3]
  PIN SEL[4]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 17.715 -2.635 18.505 -2.390 ;
      LAYER mcon ;
        RECT 18.070 -2.565 18.240 -2.395 ;
      LAYER met1 ;
        RECT 17.810 -2.770 18.430 -2.240 ;
      LAYER via ;
        RECT 18.015 -2.625 18.295 -2.345 ;
      LAYER met2 ;
        RECT 17.900 -4.360 18.370 -2.240 ;
    END
  END SEL[4]
  PIN SEL[5]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 21.075 -2.635 21.865 -2.390 ;
      LAYER mcon ;
        RECT 21.430 -2.565 21.600 -2.395 ;
      LAYER met1 ;
        RECT 21.170 -2.770 21.790 -2.240 ;
      LAYER via ;
        RECT 21.375 -2.625 21.655 -2.345 ;
      LAYER met2 ;
        RECT 21.260 -4.360 21.730 -2.240 ;
    END
  END SEL[5]
  PIN SEL[6]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 24.435 -2.635 25.225 -2.390 ;
      LAYER mcon ;
        RECT 24.790 -2.565 24.960 -2.395 ;
      LAYER met1 ;
        RECT 24.530 -2.770 25.150 -2.240 ;
      LAYER via ;
        RECT 24.735 -2.625 25.015 -2.345 ;
      LAYER met2 ;
        RECT 24.620 -4.360 25.090 -2.240 ;
    END
  END SEL[6]
  PIN SEL[7]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 27.795 -2.635 28.585 -2.390 ;
      LAYER mcon ;
        RECT 28.150 -2.565 28.320 -2.395 ;
      LAYER met1 ;
        RECT 27.890 -2.770 28.510 -2.240 ;
      LAYER via ;
        RECT 28.095 -2.625 28.375 -2.345 ;
      LAYER met2 ;
        RECT 27.980 -4.360 28.450 -2.240 ;
    END
  END SEL[7]
  PIN SEL[8]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 31.155 -2.635 31.945 -2.390 ;
      LAYER mcon ;
        RECT 31.510 -2.565 31.680 -2.395 ;
      LAYER met1 ;
        RECT 31.250 -2.770 31.870 -2.240 ;
      LAYER via ;
        RECT 31.455 -2.625 31.735 -2.345 ;
      LAYER met2 ;
        RECT 31.340 -4.360 31.810 -2.240 ;
    END
  END SEL[8]
  PIN SEL[9]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 34.515 -2.635 35.305 -2.390 ;
      LAYER mcon ;
        RECT 34.870 -2.565 35.040 -2.395 ;
      LAYER met1 ;
        RECT 34.610 -2.770 35.230 -2.240 ;
      LAYER via ;
        RECT 34.815 -2.625 35.095 -2.345 ;
      LAYER met2 ;
        RECT 34.700 -4.360 35.170 -2.240 ;
    END
  END SEL[9]
  PIN SEL[10]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 37.875 -2.635 38.665 -2.390 ;
      LAYER mcon ;
        RECT 38.230 -2.565 38.400 -2.395 ;
      LAYER met1 ;
        RECT 37.970 -2.770 38.590 -2.240 ;
      LAYER via ;
        RECT 38.175 -2.625 38.455 -2.345 ;
      LAYER met2 ;
        RECT 38.060 -4.360 38.530 -2.240 ;
    END
  END SEL[10]
  PIN SEL[11]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 41.235 -2.635 42.025 -2.390 ;
      LAYER mcon ;
        RECT 41.590 -2.565 41.760 -2.395 ;
      LAYER met1 ;
        RECT 41.330 -2.770 41.950 -2.240 ;
      LAYER via ;
        RECT 41.535 -2.625 41.815 -2.345 ;
      LAYER met2 ;
        RECT 41.420 -4.360 41.890 -2.240 ;
    END
  END SEL[11]
  PIN SEL[12]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 44.595 -2.635 45.385 -2.390 ;
      LAYER mcon ;
        RECT 44.950 -2.565 45.120 -2.395 ;
      LAYER met1 ;
        RECT 44.690 -2.770 45.310 -2.240 ;
      LAYER via ;
        RECT 44.895 -2.625 45.175 -2.345 ;
      LAYER met2 ;
        RECT 44.780 -4.360 45.250 -2.240 ;
    END
  END SEL[12]
  PIN SEL[13]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 47.955 -2.635 48.745 -2.390 ;
      LAYER mcon ;
        RECT 48.310 -2.565 48.480 -2.395 ;
      LAYER met1 ;
        RECT 48.050 -2.770 48.670 -2.240 ;
      LAYER via ;
        RECT 48.255 -2.625 48.535 -2.345 ;
      LAYER met2 ;
        RECT 48.140 -4.360 48.610 -2.240 ;
    END
  END SEL[13]
  PIN SEL[14]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 51.315 -2.635 52.105 -2.390 ;
      LAYER mcon ;
        RECT 51.670 -2.565 51.840 -2.395 ;
      LAYER met1 ;
        RECT 51.410 -2.770 52.030 -2.240 ;
      LAYER via ;
        RECT 51.615 -2.625 51.895 -2.345 ;
      LAYER met2 ;
        RECT 51.500 -4.360 51.970 -2.240 ;
    END
  END SEL[14]
  PIN SEL[15]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 54.675 -2.635 55.465 -2.390 ;
      LAYER mcon ;
        RECT 55.030 -2.565 55.200 -2.395 ;
      LAYER met1 ;
        RECT 54.770 -2.770 55.390 -2.240 ;
      LAYER via ;
        RECT 54.975 -2.625 55.255 -2.345 ;
      LAYER met2 ;
        RECT 54.860 -4.360 55.330 -2.240 ;
    END
  END SEL[15]
  PIN SEL[16]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 58.035 -2.635 58.825 -2.390 ;
      LAYER mcon ;
        RECT 58.390 -2.565 58.560 -2.395 ;
      LAYER met1 ;
        RECT 58.130 -2.770 58.750 -2.240 ;
      LAYER via ;
        RECT 58.335 -2.625 58.615 -2.345 ;
      LAYER met2 ;
        RECT 58.220 -4.360 58.690 -2.240 ;
    END
  END SEL[16]
  PIN SEL[17]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 61.395 -2.635 62.185 -2.390 ;
      LAYER mcon ;
        RECT 61.750 -2.565 61.920 -2.395 ;
      LAYER met1 ;
        RECT 61.490 -2.770 62.110 -2.240 ;
      LAYER via ;
        RECT 61.695 -2.625 61.975 -2.345 ;
      LAYER met2 ;
        RECT 61.580 -4.360 62.050 -2.240 ;
    END
  END SEL[17]
  PIN SEL[18]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 64.755 -2.635 65.545 -2.390 ;
      LAYER mcon ;
        RECT 65.110 -2.565 65.280 -2.395 ;
      LAYER met1 ;
        RECT 64.850 -2.770 65.470 -2.240 ;
      LAYER via ;
        RECT 65.055 -2.625 65.335 -2.345 ;
      LAYER met2 ;
        RECT 64.940 -4.360 65.410 -2.240 ;
    END
  END SEL[18]
  PIN SEL[19]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 68.115 -2.635 68.905 -2.390 ;
      LAYER mcon ;
        RECT 68.470 -2.565 68.640 -2.395 ;
      LAYER met1 ;
        RECT 68.210 -2.770 68.830 -2.240 ;
      LAYER via ;
        RECT 68.415 -2.625 68.695 -2.345 ;
      LAYER met2 ;
        RECT 68.300 -4.360 68.770 -2.240 ;
    END
  END SEL[19]
  PIN SEL[20]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 71.475 -2.635 72.265 -2.390 ;
      LAYER mcon ;
        RECT 71.830 -2.565 72.000 -2.395 ;
      LAYER met1 ;
        RECT 71.570 -2.770 72.190 -2.240 ;
      LAYER via ;
        RECT 71.775 -2.625 72.055 -2.345 ;
      LAYER met2 ;
        RECT 71.660 -4.360 72.130 -2.240 ;
    END
  END SEL[20]
  PIN SEL[21]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 74.835 -2.635 75.625 -2.390 ;
      LAYER mcon ;
        RECT 75.190 -2.565 75.360 -2.395 ;
      LAYER met1 ;
        RECT 74.930 -2.770 75.550 -2.240 ;
      LAYER via ;
        RECT 75.135 -2.625 75.415 -2.345 ;
      LAYER met2 ;
        RECT 75.020 -4.360 75.490 -2.240 ;
    END
  END SEL[21]
  PIN SEL[22]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 78.195 -2.635 78.985 -2.390 ;
      LAYER mcon ;
        RECT 78.550 -2.565 78.720 -2.395 ;
      LAYER met1 ;
        RECT 78.290 -2.770 78.910 -2.240 ;
      LAYER via ;
        RECT 78.495 -2.625 78.775 -2.345 ;
      LAYER met2 ;
        RECT 78.380 -4.360 78.850 -2.240 ;
    END
  END SEL[22]
  PIN SEL[23]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 81.555 -2.635 82.345 -2.390 ;
      LAYER mcon ;
        RECT 81.910 -2.565 82.080 -2.395 ;
      LAYER met1 ;
        RECT 81.650 -2.770 82.270 -2.240 ;
      LAYER via ;
        RECT 81.855 -2.625 82.135 -2.345 ;
      LAYER met2 ;
        RECT 81.740 -4.360 82.210 -2.240 ;
    END
  END SEL[23]
  PIN SEL[24]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 84.915 -2.635 85.705 -2.390 ;
      LAYER mcon ;
        RECT 85.270 -2.565 85.440 -2.395 ;
      LAYER met1 ;
        RECT 85.010 -2.770 85.630 -2.240 ;
      LAYER via ;
        RECT 85.215 -2.625 85.495 -2.345 ;
      LAYER met2 ;
        RECT 85.100 -4.360 85.570 -2.240 ;
    END
  END SEL[24]
  PIN SEL[25]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 88.275 -2.635 89.065 -2.390 ;
      LAYER mcon ;
        RECT 88.630 -2.565 88.800 -2.395 ;
      LAYER met1 ;
        RECT 88.370 -2.770 88.990 -2.240 ;
      LAYER via ;
        RECT 88.575 -2.625 88.855 -2.345 ;
      LAYER met2 ;
        RECT 88.460 -4.360 88.930 -2.240 ;
    END
  END SEL[25]
  PIN SEL[26]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 91.635 -2.635 92.425 -2.390 ;
      LAYER mcon ;
        RECT 91.990 -2.565 92.160 -2.395 ;
      LAYER met1 ;
        RECT 91.730 -2.770 92.350 -2.240 ;
      LAYER via ;
        RECT 91.935 -2.625 92.215 -2.345 ;
      LAYER met2 ;
        RECT 91.820 -4.360 92.290 -2.240 ;
    END
  END SEL[26]
  PIN SEL[27]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 94.995 -2.635 95.785 -2.390 ;
      LAYER mcon ;
        RECT 95.350 -2.565 95.520 -2.395 ;
      LAYER met1 ;
        RECT 95.090 -2.770 95.710 -2.240 ;
      LAYER via ;
        RECT 95.295 -2.625 95.575 -2.345 ;
      LAYER met2 ;
        RECT 95.180 -4.360 95.650 -2.240 ;
    END
  END SEL[27]
  PIN SEL[28]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 98.355 -2.635 99.145 -2.390 ;
      LAYER mcon ;
        RECT 98.710 -2.565 98.880 -2.395 ;
      LAYER met1 ;
        RECT 98.450 -2.770 99.070 -2.240 ;
      LAYER via ;
        RECT 98.655 -2.625 98.935 -2.345 ;
      LAYER met2 ;
        RECT 98.540 -4.360 99.010 -2.240 ;
    END
  END SEL[28]
  PIN SEL[29]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 101.715 -2.635 102.505 -2.390 ;
      LAYER mcon ;
        RECT 102.070 -2.565 102.240 -2.395 ;
      LAYER met1 ;
        RECT 101.810 -2.770 102.430 -2.240 ;
      LAYER via ;
        RECT 102.015 -2.625 102.295 -2.345 ;
      LAYER met2 ;
        RECT 101.900 -4.360 102.370 -2.240 ;
    END
  END SEL[29]
  PIN SEL[30]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 105.075 -2.635 105.865 -2.390 ;
      LAYER mcon ;
        RECT 105.430 -2.565 105.600 -2.395 ;
      LAYER met1 ;
        RECT 105.170 -2.770 105.790 -2.240 ;
      LAYER via ;
        RECT 105.375 -2.625 105.655 -2.345 ;
      LAYER met2 ;
        RECT 105.260 -4.360 105.730 -2.240 ;
    END
  END SEL[30]
  PIN SEL[31]
    ANTENNAGATEAREA 0.960000 ;
    PORT
      LAYER li1 ;
        RECT 108.435 -2.635 109.225 -2.390 ;
      LAYER mcon ;
        RECT 108.790 -2.565 108.960 -2.395 ;
      LAYER met1 ;
        RECT 108.530 -2.770 109.150 -2.240 ;
      LAYER via ;
        RECT 108.735 -2.625 109.015 -2.345 ;
      LAYER met2 ;
        RECT 108.620 -4.360 109.090 -2.240 ;
    END
  END SEL[31]
  OBS
      LAYER pwell ;
        RECT -3.490 3.785 0.130 4.215 ;
        RECT -3.340 2.585 -0.050 3.785 ;
      LAYER nwell ;
        RECT 3.430 -2.255 111.610 0.345 ;
      LAYER pwell ;
        RECT -3.340 -3.925 -0.020 -2.645 ;
        RECT 3.780 -3.925 7.100 -2.645 ;
        RECT 7.140 -3.925 10.460 -2.645 ;
        RECT 10.500 -3.925 13.820 -2.645 ;
        RECT 13.860 -3.925 17.180 -2.645 ;
        RECT 17.220 -3.925 20.540 -2.645 ;
        RECT 20.580 -3.925 23.900 -2.645 ;
        RECT 23.940 -3.925 27.260 -2.645 ;
        RECT 27.300 -3.925 30.620 -2.645 ;
        RECT 30.660 -3.925 33.980 -2.645 ;
        RECT 34.020 -3.925 37.340 -2.645 ;
        RECT 37.380 -3.925 40.700 -2.645 ;
        RECT 40.740 -3.925 44.060 -2.645 ;
        RECT 44.100 -3.925 47.420 -2.645 ;
        RECT 47.460 -3.925 50.780 -2.645 ;
        RECT 50.820 -3.925 54.140 -2.645 ;
        RECT 54.180 -3.925 57.500 -2.645 ;
        RECT 57.540 -3.925 60.860 -2.645 ;
        RECT 60.900 -3.925 64.220 -2.645 ;
        RECT 64.260 -3.925 67.580 -2.645 ;
        RECT 67.620 -3.925 70.940 -2.645 ;
        RECT 70.980 -3.925 74.300 -2.645 ;
        RECT 74.340 -3.925 77.660 -2.645 ;
        RECT 77.700 -3.925 81.020 -2.645 ;
        RECT 81.060 -3.925 84.380 -2.645 ;
        RECT 84.420 -3.925 87.740 -2.645 ;
        RECT 87.780 -3.925 91.100 -2.645 ;
        RECT 91.140 -3.925 94.460 -2.645 ;
        RECT 94.500 -3.925 97.820 -2.645 ;
        RECT 97.860 -3.925 101.180 -2.645 ;
        RECT 101.220 -3.925 104.540 -2.645 ;
        RECT 104.580 -3.925 107.900 -2.645 ;
        RECT 107.940 -3.925 111.260 -2.645 ;
        RECT -3.490 -4.355 0.130 -3.925 ;
        RECT 3.630 -4.355 111.410 -3.925 ;
      LAYER li1 ;
        RECT -3.360 3.915 0.000 4.085 ;
        RECT -2.920 3.260 -0.590 3.635 ;
        RECT -2.750 3.100 -0.590 3.260 ;
        RECT -3.270 2.575 -2.920 3.090 ;
        RECT -2.750 2.755 -1.025 3.100 ;
        RECT -3.270 2.355 -1.295 2.575 ;
        RECT -3.270 1.805 -3.015 2.355 ;
        RECT -0.410 2.120 -0.125 3.505 ;
        RECT -3.270 1.700 -2.905 1.805 ;
        RECT -3.270 0.975 -2.825 1.700 ;
        RECT -0.410 1.430 2.600 2.120 ;
        RECT -0.410 0.245 -0.125 1.430 ;
        RECT -3.185 -2.040 -2.710 -1.135 ;
        RECT -0.380 -1.190 -0.125 0.245 ;
        RECT 2.030 -1.190 2.600 1.430 ;
        RECT 3.760 -0.155 5.800 0.015 ;
        RECT 7.120 -0.155 9.160 0.015 ;
        RECT 10.480 -0.155 12.520 0.015 ;
        RECT 13.840 -0.155 15.880 0.015 ;
        RECT 17.200 -0.155 19.240 0.015 ;
        RECT 20.560 -0.155 22.600 0.015 ;
        RECT 23.920 -0.155 25.960 0.015 ;
        RECT 27.280 -0.155 29.320 0.015 ;
        RECT 30.640 -0.155 32.680 0.015 ;
        RECT 34.000 -0.155 36.040 0.015 ;
        RECT 37.360 -0.155 39.400 0.015 ;
        RECT 40.720 -0.155 42.760 0.015 ;
        RECT 44.080 -0.155 46.120 0.015 ;
        RECT 47.440 -0.155 49.480 0.015 ;
        RECT 50.800 -0.155 52.840 0.015 ;
        RECT 54.160 -0.155 56.200 0.015 ;
        RECT 57.520 -0.155 59.560 0.015 ;
        RECT 60.880 -0.155 62.920 0.015 ;
        RECT 64.240 -0.155 66.280 0.015 ;
        RECT 67.600 -0.155 69.640 0.015 ;
        RECT 70.960 -0.155 73.000 0.015 ;
        RECT 74.320 -0.155 76.360 0.015 ;
        RECT 77.680 -0.155 79.720 0.015 ;
        RECT 81.040 -0.155 83.080 0.015 ;
        RECT 84.400 -0.155 86.440 0.015 ;
        RECT 87.760 -0.155 89.800 0.015 ;
        RECT 91.120 -0.155 93.160 0.015 ;
        RECT 94.480 -0.155 96.520 0.015 ;
        RECT 97.840 -0.155 99.880 0.015 ;
        RECT 101.200 -0.155 103.240 0.015 ;
        RECT 104.560 -0.155 106.600 0.015 ;
        RECT 107.920 -0.155 109.960 0.015 ;
        RECT -0.380 -1.850 2.600 -1.190 ;
        RECT -0.380 -2.015 -0.125 -1.850 ;
        RECT -3.185 -2.210 -1.295 -2.040 ;
        RECT -3.185 -2.805 -3.015 -2.210 ;
        RECT -1.885 -2.415 -1.295 -2.210 ;
        RECT -0.325 -2.685 -0.125 -2.015 ;
        RECT -3.185 -3.235 -2.980 -2.805 ;
        RECT -2.810 -3.150 -1.085 -2.805 ;
        RECT -2.810 -3.405 -0.560 -3.150 ;
        RECT -2.890 -3.775 -0.560 -3.405 ;
        RECT -0.380 -3.565 -0.125 -2.685 ;
        RECT 3.935 -2.040 4.410 -1.135 ;
        RECT 4.590 -1.430 6.560 -0.385 ;
        RECT 4.590 -1.860 6.035 -1.430 ;
        RECT 7.295 -2.040 7.770 -1.135 ;
        RECT 7.950 -1.430 9.920 -0.385 ;
        RECT 7.950 -1.860 9.395 -1.430 ;
        RECT 10.655 -2.040 11.130 -1.135 ;
        RECT 11.310 -1.430 13.280 -0.385 ;
        RECT 11.310 -1.860 12.755 -1.430 ;
        RECT 14.015 -2.040 14.490 -1.135 ;
        RECT 14.670 -1.430 16.640 -0.385 ;
        RECT 14.670 -1.860 16.115 -1.430 ;
        RECT 17.375 -2.040 17.850 -1.135 ;
        RECT 18.030 -1.430 20.000 -0.385 ;
        RECT 18.030 -1.860 19.475 -1.430 ;
        RECT 20.735 -2.040 21.210 -1.135 ;
        RECT 21.390 -1.430 23.360 -0.385 ;
        RECT 21.390 -1.860 22.835 -1.430 ;
        RECT 24.095 -2.040 24.570 -1.135 ;
        RECT 24.750 -1.430 26.720 -0.385 ;
        RECT 24.750 -1.860 26.195 -1.430 ;
        RECT 27.455 -2.040 27.930 -1.135 ;
        RECT 28.110 -1.430 30.080 -0.385 ;
        RECT 28.110 -1.860 29.555 -1.430 ;
        RECT 30.815 -2.040 31.290 -1.135 ;
        RECT 31.470 -1.430 33.440 -0.385 ;
        RECT 31.470 -1.860 32.915 -1.430 ;
        RECT 34.175 -2.040 34.650 -1.135 ;
        RECT 34.830 -1.430 36.800 -0.385 ;
        RECT 34.830 -1.860 36.275 -1.430 ;
        RECT 37.535 -2.040 38.010 -1.135 ;
        RECT 38.190 -1.430 40.160 -0.385 ;
        RECT 38.190 -1.860 39.635 -1.430 ;
        RECT 40.895 -2.040 41.370 -1.135 ;
        RECT 41.550 -1.430 43.520 -0.385 ;
        RECT 41.550 -1.860 42.995 -1.430 ;
        RECT 44.255 -2.040 44.730 -1.135 ;
        RECT 44.910 -1.430 46.880 -0.385 ;
        RECT 44.910 -1.860 46.355 -1.430 ;
        RECT 47.615 -2.040 48.090 -1.135 ;
        RECT 48.270 -1.430 50.240 -0.385 ;
        RECT 48.270 -1.860 49.715 -1.430 ;
        RECT 50.975 -2.040 51.450 -1.135 ;
        RECT 51.630 -1.430 53.600 -0.385 ;
        RECT 51.630 -1.860 53.075 -1.430 ;
        RECT 54.335 -2.040 54.810 -1.135 ;
        RECT 54.990 -1.430 56.960 -0.385 ;
        RECT 54.990 -1.860 56.435 -1.430 ;
        RECT 57.695 -2.040 58.170 -1.135 ;
        RECT 58.350 -1.430 60.320 -0.385 ;
        RECT 58.350 -1.860 59.795 -1.430 ;
        RECT 61.055 -2.040 61.530 -1.135 ;
        RECT 61.710 -1.430 63.680 -0.385 ;
        RECT 61.710 -1.860 63.155 -1.430 ;
        RECT 64.415 -2.040 64.890 -1.135 ;
        RECT 65.070 -1.430 67.040 -0.385 ;
        RECT 65.070 -1.860 66.515 -1.430 ;
        RECT 67.775 -2.040 68.250 -1.135 ;
        RECT 68.430 -1.430 70.400 -0.385 ;
        RECT 68.430 -1.860 69.875 -1.430 ;
        RECT 71.135 -2.040 71.610 -1.135 ;
        RECT 71.790 -1.430 73.760 -0.385 ;
        RECT 71.790 -1.860 73.235 -1.430 ;
        RECT 74.495 -2.040 74.970 -1.135 ;
        RECT 75.150 -1.430 77.120 -0.385 ;
        RECT 75.150 -1.860 76.595 -1.430 ;
        RECT 77.855 -2.040 78.330 -1.135 ;
        RECT 78.510 -1.430 80.480 -0.385 ;
        RECT 78.510 -1.860 79.955 -1.430 ;
        RECT 81.215 -2.040 81.690 -1.135 ;
        RECT 81.870 -1.430 83.840 -0.385 ;
        RECT 81.870 -1.860 83.315 -1.430 ;
        RECT 84.575 -2.040 85.050 -1.135 ;
        RECT 85.230 -1.430 87.200 -0.385 ;
        RECT 85.230 -1.860 86.675 -1.430 ;
        RECT 87.935 -2.040 88.410 -1.135 ;
        RECT 88.590 -1.430 90.560 -0.385 ;
        RECT 88.590 -1.860 90.035 -1.430 ;
        RECT 91.295 -2.040 91.770 -1.135 ;
        RECT 91.950 -1.430 93.920 -0.385 ;
        RECT 91.950 -1.860 93.395 -1.430 ;
        RECT 94.655 -2.040 95.130 -1.135 ;
        RECT 95.310 -1.430 97.280 -0.385 ;
        RECT 95.310 -1.860 96.755 -1.430 ;
        RECT 98.015 -2.040 98.490 -1.135 ;
        RECT 98.670 -1.430 100.640 -0.385 ;
        RECT 98.670 -1.860 100.115 -1.430 ;
        RECT 101.375 -2.040 101.850 -1.135 ;
        RECT 102.030 -1.430 104.000 -0.385 ;
        RECT 102.030 -1.860 103.475 -1.430 ;
        RECT 104.735 -2.040 105.210 -1.135 ;
        RECT 105.390 -1.430 107.360 -0.385 ;
        RECT 105.390 -1.860 106.835 -1.430 ;
        RECT 108.095 -2.040 108.570 -1.135 ;
        RECT 108.750 -1.430 110.720 -0.385 ;
        RECT 108.750 -1.860 110.195 -1.430 ;
        RECT 3.935 -2.210 5.825 -2.040 ;
        RECT 3.935 -2.805 4.105 -2.210 ;
        RECT 5.235 -2.415 5.825 -2.210 ;
        RECT 7.295 -2.210 9.185 -2.040 ;
        RECT 7.295 -2.805 7.465 -2.210 ;
        RECT 8.595 -2.415 9.185 -2.210 ;
        RECT 10.655 -2.210 12.545 -2.040 ;
        RECT 10.655 -2.805 10.825 -2.210 ;
        RECT 11.955 -2.415 12.545 -2.210 ;
        RECT 14.015 -2.210 15.905 -2.040 ;
        RECT 14.015 -2.805 14.185 -2.210 ;
        RECT 15.315 -2.415 15.905 -2.210 ;
        RECT 17.375 -2.210 19.265 -2.040 ;
        RECT 17.375 -2.805 17.545 -2.210 ;
        RECT 18.675 -2.415 19.265 -2.210 ;
        RECT 20.735 -2.210 22.625 -2.040 ;
        RECT 20.735 -2.805 20.905 -2.210 ;
        RECT 22.035 -2.415 22.625 -2.210 ;
        RECT 24.095 -2.210 25.985 -2.040 ;
        RECT 24.095 -2.805 24.265 -2.210 ;
        RECT 25.395 -2.415 25.985 -2.210 ;
        RECT 27.455 -2.210 29.345 -2.040 ;
        RECT 27.455 -2.805 27.625 -2.210 ;
        RECT 28.755 -2.415 29.345 -2.210 ;
        RECT 30.815 -2.210 32.705 -2.040 ;
        RECT 30.815 -2.805 30.985 -2.210 ;
        RECT 32.115 -2.415 32.705 -2.210 ;
        RECT 34.175 -2.210 36.065 -2.040 ;
        RECT 34.175 -2.805 34.345 -2.210 ;
        RECT 35.475 -2.415 36.065 -2.210 ;
        RECT 37.535 -2.210 39.425 -2.040 ;
        RECT 37.535 -2.805 37.705 -2.210 ;
        RECT 38.835 -2.415 39.425 -2.210 ;
        RECT 40.895 -2.210 42.785 -2.040 ;
        RECT 40.895 -2.805 41.065 -2.210 ;
        RECT 42.195 -2.415 42.785 -2.210 ;
        RECT 44.255 -2.210 46.145 -2.040 ;
        RECT 44.255 -2.805 44.425 -2.210 ;
        RECT 45.555 -2.415 46.145 -2.210 ;
        RECT 47.615 -2.210 49.505 -2.040 ;
        RECT 47.615 -2.805 47.785 -2.210 ;
        RECT 48.915 -2.415 49.505 -2.210 ;
        RECT 50.975 -2.210 52.865 -2.040 ;
        RECT 50.975 -2.805 51.145 -2.210 ;
        RECT 52.275 -2.415 52.865 -2.210 ;
        RECT 54.335 -2.210 56.225 -2.040 ;
        RECT 54.335 -2.805 54.505 -2.210 ;
        RECT 55.635 -2.415 56.225 -2.210 ;
        RECT 57.695 -2.210 59.585 -2.040 ;
        RECT 57.695 -2.805 57.865 -2.210 ;
        RECT 58.995 -2.415 59.585 -2.210 ;
        RECT 61.055 -2.210 62.945 -2.040 ;
        RECT 61.055 -2.805 61.225 -2.210 ;
        RECT 62.355 -2.415 62.945 -2.210 ;
        RECT 64.415 -2.210 66.305 -2.040 ;
        RECT 64.415 -2.805 64.585 -2.210 ;
        RECT 65.715 -2.415 66.305 -2.210 ;
        RECT 67.775 -2.210 69.665 -2.040 ;
        RECT 67.775 -2.805 67.945 -2.210 ;
        RECT 69.075 -2.415 69.665 -2.210 ;
        RECT 71.135 -2.210 73.025 -2.040 ;
        RECT 71.135 -2.805 71.305 -2.210 ;
        RECT 72.435 -2.415 73.025 -2.210 ;
        RECT 74.495 -2.210 76.385 -2.040 ;
        RECT 74.495 -2.805 74.665 -2.210 ;
        RECT 75.795 -2.415 76.385 -2.210 ;
        RECT 77.855 -2.210 79.745 -2.040 ;
        RECT 77.855 -2.805 78.025 -2.210 ;
        RECT 79.155 -2.415 79.745 -2.210 ;
        RECT 81.215 -2.210 83.105 -2.040 ;
        RECT 81.215 -2.805 81.385 -2.210 ;
        RECT 82.515 -2.415 83.105 -2.210 ;
        RECT 84.575 -2.210 86.465 -2.040 ;
        RECT 84.575 -2.805 84.745 -2.210 ;
        RECT 85.875 -2.415 86.465 -2.210 ;
        RECT 87.935 -2.210 89.825 -2.040 ;
        RECT 87.935 -2.805 88.105 -2.210 ;
        RECT 89.235 -2.415 89.825 -2.210 ;
        RECT 91.295 -2.210 93.185 -2.040 ;
        RECT 91.295 -2.805 91.465 -2.210 ;
        RECT 92.595 -2.415 93.185 -2.210 ;
        RECT 94.655 -2.210 96.545 -2.040 ;
        RECT 94.655 -2.805 94.825 -2.210 ;
        RECT 95.955 -2.415 96.545 -2.210 ;
        RECT 98.015 -2.210 99.905 -2.040 ;
        RECT 98.015 -2.805 98.185 -2.210 ;
        RECT 99.315 -2.415 99.905 -2.210 ;
        RECT 101.375 -2.210 103.265 -2.040 ;
        RECT 101.375 -2.805 101.545 -2.210 ;
        RECT 102.675 -2.415 103.265 -2.210 ;
        RECT 104.735 -2.210 106.625 -2.040 ;
        RECT 104.735 -2.805 104.905 -2.210 ;
        RECT 106.035 -2.415 106.625 -2.210 ;
        RECT 108.095 -2.210 109.985 -2.040 ;
        RECT 108.095 -2.805 108.265 -2.210 ;
        RECT 109.395 -2.415 109.985 -2.210 ;
        RECT 3.935 -3.235 4.140 -2.805 ;
        RECT 4.310 -3.150 6.035 -2.805 ;
        RECT 4.310 -3.405 6.560 -3.150 ;
        RECT 7.295 -3.235 7.500 -2.805 ;
        RECT 7.670 -3.150 9.395 -2.805 ;
        RECT 7.670 -3.405 9.920 -3.150 ;
        RECT 10.655 -3.235 10.860 -2.805 ;
        RECT 11.030 -3.150 12.755 -2.805 ;
        RECT 11.030 -3.405 13.280 -3.150 ;
        RECT 14.015 -3.235 14.220 -2.805 ;
        RECT 14.390 -3.150 16.115 -2.805 ;
        RECT 14.390 -3.405 16.640 -3.150 ;
        RECT 17.375 -3.235 17.580 -2.805 ;
        RECT 17.750 -3.150 19.475 -2.805 ;
        RECT 17.750 -3.405 20.000 -3.150 ;
        RECT 20.735 -3.235 20.940 -2.805 ;
        RECT 21.110 -3.150 22.835 -2.805 ;
        RECT 21.110 -3.405 23.360 -3.150 ;
        RECT 24.095 -3.235 24.300 -2.805 ;
        RECT 24.470 -3.150 26.195 -2.805 ;
        RECT 24.470 -3.405 26.720 -3.150 ;
        RECT 27.455 -3.235 27.660 -2.805 ;
        RECT 27.830 -3.150 29.555 -2.805 ;
        RECT 27.830 -3.405 30.080 -3.150 ;
        RECT 30.815 -3.235 31.020 -2.805 ;
        RECT 31.190 -3.150 32.915 -2.805 ;
        RECT 31.190 -3.405 33.440 -3.150 ;
        RECT 34.175 -3.235 34.380 -2.805 ;
        RECT 34.550 -3.150 36.275 -2.805 ;
        RECT 34.550 -3.405 36.800 -3.150 ;
        RECT 37.535 -3.235 37.740 -2.805 ;
        RECT 37.910 -3.150 39.635 -2.805 ;
        RECT 37.910 -3.405 40.160 -3.150 ;
        RECT 40.895 -3.235 41.100 -2.805 ;
        RECT 41.270 -3.150 42.995 -2.805 ;
        RECT 41.270 -3.405 43.520 -3.150 ;
        RECT 44.255 -3.235 44.460 -2.805 ;
        RECT 44.630 -3.150 46.355 -2.805 ;
        RECT 44.630 -3.405 46.880 -3.150 ;
        RECT 47.615 -3.235 47.820 -2.805 ;
        RECT 47.990 -3.150 49.715 -2.805 ;
        RECT 47.990 -3.405 50.240 -3.150 ;
        RECT 50.975 -3.235 51.180 -2.805 ;
        RECT 51.350 -3.150 53.075 -2.805 ;
        RECT 51.350 -3.405 53.600 -3.150 ;
        RECT 54.335 -3.235 54.540 -2.805 ;
        RECT 54.710 -3.150 56.435 -2.805 ;
        RECT 54.710 -3.405 56.960 -3.150 ;
        RECT 57.695 -3.235 57.900 -2.805 ;
        RECT 58.070 -3.150 59.795 -2.805 ;
        RECT 58.070 -3.405 60.320 -3.150 ;
        RECT 61.055 -3.235 61.260 -2.805 ;
        RECT 61.430 -3.150 63.155 -2.805 ;
        RECT 61.430 -3.405 63.680 -3.150 ;
        RECT 64.415 -3.235 64.620 -2.805 ;
        RECT 64.790 -3.150 66.515 -2.805 ;
        RECT 64.790 -3.405 67.040 -3.150 ;
        RECT 67.775 -3.235 67.980 -2.805 ;
        RECT 68.150 -3.150 69.875 -2.805 ;
        RECT 68.150 -3.405 70.400 -3.150 ;
        RECT 71.135 -3.235 71.340 -2.805 ;
        RECT 71.510 -3.150 73.235 -2.805 ;
        RECT 71.510 -3.405 73.760 -3.150 ;
        RECT 74.495 -3.235 74.700 -2.805 ;
        RECT 74.870 -3.150 76.595 -2.805 ;
        RECT 74.870 -3.405 77.120 -3.150 ;
        RECT 77.855 -3.235 78.060 -2.805 ;
        RECT 78.230 -3.150 79.955 -2.805 ;
        RECT 78.230 -3.405 80.480 -3.150 ;
        RECT 81.215 -3.235 81.420 -2.805 ;
        RECT 81.590 -3.150 83.315 -2.805 ;
        RECT 81.590 -3.405 83.840 -3.150 ;
        RECT 84.575 -3.235 84.780 -2.805 ;
        RECT 84.950 -3.150 86.675 -2.805 ;
        RECT 84.950 -3.405 87.200 -3.150 ;
        RECT 87.935 -3.235 88.140 -2.805 ;
        RECT 88.310 -3.150 90.035 -2.805 ;
        RECT 88.310 -3.405 90.560 -3.150 ;
        RECT 91.295 -3.235 91.500 -2.805 ;
        RECT 91.670 -3.150 93.395 -2.805 ;
        RECT 91.670 -3.405 93.920 -3.150 ;
        RECT 94.655 -3.235 94.860 -2.805 ;
        RECT 95.030 -3.150 96.755 -2.805 ;
        RECT 95.030 -3.405 97.280 -3.150 ;
        RECT 98.015 -3.235 98.220 -2.805 ;
        RECT 98.390 -3.150 100.115 -2.805 ;
        RECT 98.390 -3.405 100.640 -3.150 ;
        RECT 101.375 -3.235 101.580 -2.805 ;
        RECT 101.750 -3.150 103.475 -2.805 ;
        RECT 101.750 -3.405 104.000 -3.150 ;
        RECT 104.735 -3.235 104.940 -2.805 ;
        RECT 105.110 -3.150 106.835 -2.805 ;
        RECT 105.110 -3.405 107.360 -3.150 ;
        RECT 108.095 -3.235 108.300 -2.805 ;
        RECT 108.470 -3.150 110.195 -2.805 ;
        RECT 108.470 -3.405 110.720 -3.150 ;
        RECT 4.230 -3.775 6.560 -3.405 ;
        RECT 7.590 -3.775 9.920 -3.405 ;
        RECT 10.950 -3.775 13.280 -3.405 ;
        RECT 14.310 -3.775 16.640 -3.405 ;
        RECT 17.670 -3.775 20.000 -3.405 ;
        RECT 21.030 -3.775 23.360 -3.405 ;
        RECT 24.390 -3.775 26.720 -3.405 ;
        RECT 27.750 -3.775 30.080 -3.405 ;
        RECT 31.110 -3.775 33.440 -3.405 ;
        RECT 34.470 -3.775 36.800 -3.405 ;
        RECT 37.830 -3.775 40.160 -3.405 ;
        RECT 41.190 -3.775 43.520 -3.405 ;
        RECT 44.550 -3.775 46.880 -3.405 ;
        RECT 47.910 -3.775 50.240 -3.405 ;
        RECT 51.270 -3.775 53.600 -3.405 ;
        RECT 54.630 -3.775 56.960 -3.405 ;
        RECT 57.990 -3.775 60.320 -3.405 ;
        RECT 61.350 -3.775 63.680 -3.405 ;
        RECT 64.710 -3.775 67.040 -3.405 ;
        RECT 68.070 -3.775 70.400 -3.405 ;
        RECT 71.430 -3.775 73.760 -3.405 ;
        RECT 74.790 -3.775 77.120 -3.405 ;
        RECT 78.150 -3.775 80.480 -3.405 ;
        RECT 81.510 -3.775 83.840 -3.405 ;
        RECT 84.870 -3.775 87.200 -3.405 ;
        RECT 88.230 -3.775 90.560 -3.405 ;
        RECT 91.590 -3.775 93.920 -3.405 ;
        RECT 94.950 -3.775 97.280 -3.405 ;
        RECT 98.310 -3.775 100.640 -3.405 ;
        RECT 101.670 -3.775 104.000 -3.405 ;
        RECT 105.030 -3.775 107.360 -3.405 ;
        RECT 108.390 -3.775 110.720 -3.405 ;
        RECT -3.360 -4.225 0.000 -4.055 ;
        RECT 3.760 -4.225 111.280 -4.055 ;
      LAYER mcon ;
        RECT -3.205 3.915 -3.035 4.085 ;
        RECT -2.725 3.915 -2.555 4.085 ;
        RECT -2.245 3.915 -2.075 4.085 ;
        RECT -1.765 3.915 -1.595 4.085 ;
        RECT -1.285 3.915 -1.115 4.085 ;
        RECT -0.805 3.915 -0.635 4.085 ;
        RECT -0.325 3.915 -0.155 4.085 ;
        RECT -2.920 3.435 -2.750 3.605 ;
        RECT -2.560 3.435 -2.390 3.605 ;
        RECT -2.200 3.435 -2.030 3.605 ;
        RECT -1.840 3.435 -1.670 3.605 ;
        RECT -1.480 3.435 -1.310 3.605 ;
        RECT -1.120 3.435 -0.950 3.605 ;
        RECT -0.760 3.435 -0.590 3.605 ;
        RECT 2.230 -0.235 2.400 -0.065 ;
        RECT 3.915 -0.155 4.085 0.015 ;
        RECT 4.395 -0.155 4.565 0.015 ;
        RECT 4.875 -0.155 5.045 0.015 ;
        RECT 5.355 -0.155 5.525 0.015 ;
        RECT 7.275 -0.155 7.445 0.015 ;
        RECT 7.755 -0.155 7.925 0.015 ;
        RECT 8.235 -0.155 8.405 0.015 ;
        RECT 8.715 -0.155 8.885 0.015 ;
        RECT 10.635 -0.155 10.805 0.015 ;
        RECT 11.115 -0.155 11.285 0.015 ;
        RECT 11.595 -0.155 11.765 0.015 ;
        RECT 12.075 -0.155 12.245 0.015 ;
        RECT 13.995 -0.155 14.165 0.015 ;
        RECT 14.475 -0.155 14.645 0.015 ;
        RECT 14.955 -0.155 15.125 0.015 ;
        RECT 15.435 -0.155 15.605 0.015 ;
        RECT 17.355 -0.155 17.525 0.015 ;
        RECT 17.835 -0.155 18.005 0.015 ;
        RECT 18.315 -0.155 18.485 0.015 ;
        RECT 18.795 -0.155 18.965 0.015 ;
        RECT 20.715 -0.155 20.885 0.015 ;
        RECT 21.195 -0.155 21.365 0.015 ;
        RECT 21.675 -0.155 21.845 0.015 ;
        RECT 22.155 -0.155 22.325 0.015 ;
        RECT 24.075 -0.155 24.245 0.015 ;
        RECT 24.555 -0.155 24.725 0.015 ;
        RECT 25.035 -0.155 25.205 0.015 ;
        RECT 25.515 -0.155 25.685 0.015 ;
        RECT 27.435 -0.155 27.605 0.015 ;
        RECT 27.915 -0.155 28.085 0.015 ;
        RECT 28.395 -0.155 28.565 0.015 ;
        RECT 28.875 -0.155 29.045 0.015 ;
        RECT 30.795 -0.155 30.965 0.015 ;
        RECT 31.275 -0.155 31.445 0.015 ;
        RECT 31.755 -0.155 31.925 0.015 ;
        RECT 32.235 -0.155 32.405 0.015 ;
        RECT 34.155 -0.155 34.325 0.015 ;
        RECT 34.635 -0.155 34.805 0.015 ;
        RECT 35.115 -0.155 35.285 0.015 ;
        RECT 35.595 -0.155 35.765 0.015 ;
        RECT 37.515 -0.155 37.685 0.015 ;
        RECT 37.995 -0.155 38.165 0.015 ;
        RECT 38.475 -0.155 38.645 0.015 ;
        RECT 38.955 -0.155 39.125 0.015 ;
        RECT 40.875 -0.155 41.045 0.015 ;
        RECT 41.355 -0.155 41.525 0.015 ;
        RECT 41.835 -0.155 42.005 0.015 ;
        RECT 42.315 -0.155 42.485 0.015 ;
        RECT 44.235 -0.155 44.405 0.015 ;
        RECT 44.715 -0.155 44.885 0.015 ;
        RECT 45.195 -0.155 45.365 0.015 ;
        RECT 45.675 -0.155 45.845 0.015 ;
        RECT 47.595 -0.155 47.765 0.015 ;
        RECT 48.075 -0.155 48.245 0.015 ;
        RECT 48.555 -0.155 48.725 0.015 ;
        RECT 49.035 -0.155 49.205 0.015 ;
        RECT 50.955 -0.155 51.125 0.015 ;
        RECT 51.435 -0.155 51.605 0.015 ;
        RECT 51.915 -0.155 52.085 0.015 ;
        RECT 52.395 -0.155 52.565 0.015 ;
        RECT 54.315 -0.155 54.485 0.015 ;
        RECT 54.795 -0.155 54.965 0.015 ;
        RECT 55.275 -0.155 55.445 0.015 ;
        RECT 55.755 -0.155 55.925 0.015 ;
        RECT 57.675 -0.155 57.845 0.015 ;
        RECT 58.155 -0.155 58.325 0.015 ;
        RECT 58.635 -0.155 58.805 0.015 ;
        RECT 59.115 -0.155 59.285 0.015 ;
        RECT 61.035 -0.155 61.205 0.015 ;
        RECT 61.515 -0.155 61.685 0.015 ;
        RECT 61.995 -0.155 62.165 0.015 ;
        RECT 62.475 -0.155 62.645 0.015 ;
        RECT 64.395 -0.155 64.565 0.015 ;
        RECT 64.875 -0.155 65.045 0.015 ;
        RECT 65.355 -0.155 65.525 0.015 ;
        RECT 65.835 -0.155 66.005 0.015 ;
        RECT 67.755 -0.155 67.925 0.015 ;
        RECT 68.235 -0.155 68.405 0.015 ;
        RECT 68.715 -0.155 68.885 0.015 ;
        RECT 69.195 -0.155 69.365 0.015 ;
        RECT 71.115 -0.155 71.285 0.015 ;
        RECT 71.595 -0.155 71.765 0.015 ;
        RECT 72.075 -0.155 72.245 0.015 ;
        RECT 72.555 -0.155 72.725 0.015 ;
        RECT 74.475 -0.155 74.645 0.015 ;
        RECT 74.955 -0.155 75.125 0.015 ;
        RECT 75.435 -0.155 75.605 0.015 ;
        RECT 75.915 -0.155 76.085 0.015 ;
        RECT 77.835 -0.155 78.005 0.015 ;
        RECT 78.315 -0.155 78.485 0.015 ;
        RECT 78.795 -0.155 78.965 0.015 ;
        RECT 79.275 -0.155 79.445 0.015 ;
        RECT 81.195 -0.155 81.365 0.015 ;
        RECT 81.675 -0.155 81.845 0.015 ;
        RECT 82.155 -0.155 82.325 0.015 ;
        RECT 82.635 -0.155 82.805 0.015 ;
        RECT 84.555 -0.155 84.725 0.015 ;
        RECT 85.035 -0.155 85.205 0.015 ;
        RECT 85.515 -0.155 85.685 0.015 ;
        RECT 85.995 -0.155 86.165 0.015 ;
        RECT 87.915 -0.155 88.085 0.015 ;
        RECT 88.395 -0.155 88.565 0.015 ;
        RECT 88.875 -0.155 89.045 0.015 ;
        RECT 89.355 -0.155 89.525 0.015 ;
        RECT 91.275 -0.155 91.445 0.015 ;
        RECT 91.755 -0.155 91.925 0.015 ;
        RECT 92.235 -0.155 92.405 0.015 ;
        RECT 92.715 -0.155 92.885 0.015 ;
        RECT 94.635 -0.155 94.805 0.015 ;
        RECT 95.115 -0.155 95.285 0.015 ;
        RECT 95.595 -0.155 95.765 0.015 ;
        RECT 96.075 -0.155 96.245 0.015 ;
        RECT 97.995 -0.155 98.165 0.015 ;
        RECT 98.475 -0.155 98.645 0.015 ;
        RECT 98.955 -0.155 99.125 0.015 ;
        RECT 99.435 -0.155 99.605 0.015 ;
        RECT 101.355 -0.155 101.525 0.015 ;
        RECT 101.835 -0.155 102.005 0.015 ;
        RECT 102.315 -0.155 102.485 0.015 ;
        RECT 102.795 -0.155 102.965 0.015 ;
        RECT 104.715 -0.155 104.885 0.015 ;
        RECT 105.195 -0.155 105.365 0.015 ;
        RECT 105.675 -0.155 105.845 0.015 ;
        RECT 106.155 -0.155 106.325 0.015 ;
        RECT 108.075 -0.155 108.245 0.015 ;
        RECT 108.555 -0.155 108.725 0.015 ;
        RECT 109.035 -0.155 109.205 0.015 ;
        RECT 109.515 -0.155 109.685 0.015 ;
        RECT 2.230 -0.595 2.400 -0.425 ;
        RECT 4.590 -0.635 4.760 -0.465 ;
        RECT 4.950 -0.635 5.120 -0.465 ;
        RECT 5.310 -0.635 5.480 -0.465 ;
        RECT 5.670 -0.635 5.840 -0.465 ;
        RECT 6.030 -0.635 6.200 -0.465 ;
        RECT 6.390 -0.635 6.560 -0.465 ;
        RECT 7.950 -0.635 8.120 -0.465 ;
        RECT 8.310 -0.635 8.480 -0.465 ;
        RECT 8.670 -0.635 8.840 -0.465 ;
        RECT 9.030 -0.635 9.200 -0.465 ;
        RECT 9.390 -0.635 9.560 -0.465 ;
        RECT 9.750 -0.635 9.920 -0.465 ;
        RECT 11.310 -0.635 11.480 -0.465 ;
        RECT 11.670 -0.635 11.840 -0.465 ;
        RECT 12.030 -0.635 12.200 -0.465 ;
        RECT 12.390 -0.635 12.560 -0.465 ;
        RECT 12.750 -0.635 12.920 -0.465 ;
        RECT 13.110 -0.635 13.280 -0.465 ;
        RECT 14.670 -0.635 14.840 -0.465 ;
        RECT 15.030 -0.635 15.200 -0.465 ;
        RECT 15.390 -0.635 15.560 -0.465 ;
        RECT 15.750 -0.635 15.920 -0.465 ;
        RECT 16.110 -0.635 16.280 -0.465 ;
        RECT 16.470 -0.635 16.640 -0.465 ;
        RECT 18.030 -0.635 18.200 -0.465 ;
        RECT 18.390 -0.635 18.560 -0.465 ;
        RECT 18.750 -0.635 18.920 -0.465 ;
        RECT 19.110 -0.635 19.280 -0.465 ;
        RECT 19.470 -0.635 19.640 -0.465 ;
        RECT 19.830 -0.635 20.000 -0.465 ;
        RECT 21.390 -0.635 21.560 -0.465 ;
        RECT 21.750 -0.635 21.920 -0.465 ;
        RECT 22.110 -0.635 22.280 -0.465 ;
        RECT 22.470 -0.635 22.640 -0.465 ;
        RECT 22.830 -0.635 23.000 -0.465 ;
        RECT 23.190 -0.635 23.360 -0.465 ;
        RECT 24.750 -0.635 24.920 -0.465 ;
        RECT 25.110 -0.635 25.280 -0.465 ;
        RECT 25.470 -0.635 25.640 -0.465 ;
        RECT 25.830 -0.635 26.000 -0.465 ;
        RECT 26.190 -0.635 26.360 -0.465 ;
        RECT 26.550 -0.635 26.720 -0.465 ;
        RECT 28.110 -0.635 28.280 -0.465 ;
        RECT 28.470 -0.635 28.640 -0.465 ;
        RECT 28.830 -0.635 29.000 -0.465 ;
        RECT 29.190 -0.635 29.360 -0.465 ;
        RECT 29.550 -0.635 29.720 -0.465 ;
        RECT 29.910 -0.635 30.080 -0.465 ;
        RECT 31.470 -0.635 31.640 -0.465 ;
        RECT 31.830 -0.635 32.000 -0.465 ;
        RECT 32.190 -0.635 32.360 -0.465 ;
        RECT 32.550 -0.635 32.720 -0.465 ;
        RECT 32.910 -0.635 33.080 -0.465 ;
        RECT 33.270 -0.635 33.440 -0.465 ;
        RECT 34.830 -0.635 35.000 -0.465 ;
        RECT 35.190 -0.635 35.360 -0.465 ;
        RECT 35.550 -0.635 35.720 -0.465 ;
        RECT 35.910 -0.635 36.080 -0.465 ;
        RECT 36.270 -0.635 36.440 -0.465 ;
        RECT 36.630 -0.635 36.800 -0.465 ;
        RECT 38.190 -0.635 38.360 -0.465 ;
        RECT 38.550 -0.635 38.720 -0.465 ;
        RECT 38.910 -0.635 39.080 -0.465 ;
        RECT 39.270 -0.635 39.440 -0.465 ;
        RECT 39.630 -0.635 39.800 -0.465 ;
        RECT 39.990 -0.635 40.160 -0.465 ;
        RECT 41.550 -0.635 41.720 -0.465 ;
        RECT 41.910 -0.635 42.080 -0.465 ;
        RECT 42.270 -0.635 42.440 -0.465 ;
        RECT 42.630 -0.635 42.800 -0.465 ;
        RECT 42.990 -0.635 43.160 -0.465 ;
        RECT 43.350 -0.635 43.520 -0.465 ;
        RECT 44.910 -0.635 45.080 -0.465 ;
        RECT 45.270 -0.635 45.440 -0.465 ;
        RECT 45.630 -0.635 45.800 -0.465 ;
        RECT 45.990 -0.635 46.160 -0.465 ;
        RECT 46.350 -0.635 46.520 -0.465 ;
        RECT 46.710 -0.635 46.880 -0.465 ;
        RECT 48.270 -0.635 48.440 -0.465 ;
        RECT 48.630 -0.635 48.800 -0.465 ;
        RECT 48.990 -0.635 49.160 -0.465 ;
        RECT 49.350 -0.635 49.520 -0.465 ;
        RECT 49.710 -0.635 49.880 -0.465 ;
        RECT 50.070 -0.635 50.240 -0.465 ;
        RECT 51.630 -0.635 51.800 -0.465 ;
        RECT 51.990 -0.635 52.160 -0.465 ;
        RECT 52.350 -0.635 52.520 -0.465 ;
        RECT 52.710 -0.635 52.880 -0.465 ;
        RECT 53.070 -0.635 53.240 -0.465 ;
        RECT 53.430 -0.635 53.600 -0.465 ;
        RECT 54.990 -0.635 55.160 -0.465 ;
        RECT 55.350 -0.635 55.520 -0.465 ;
        RECT 55.710 -0.635 55.880 -0.465 ;
        RECT 56.070 -0.635 56.240 -0.465 ;
        RECT 56.430 -0.635 56.600 -0.465 ;
        RECT 56.790 -0.635 56.960 -0.465 ;
        RECT 58.350 -0.635 58.520 -0.465 ;
        RECT 58.710 -0.635 58.880 -0.465 ;
        RECT 59.070 -0.635 59.240 -0.465 ;
        RECT 59.430 -0.635 59.600 -0.465 ;
        RECT 59.790 -0.635 59.960 -0.465 ;
        RECT 60.150 -0.635 60.320 -0.465 ;
        RECT 61.710 -0.635 61.880 -0.465 ;
        RECT 62.070 -0.635 62.240 -0.465 ;
        RECT 62.430 -0.635 62.600 -0.465 ;
        RECT 62.790 -0.635 62.960 -0.465 ;
        RECT 63.150 -0.635 63.320 -0.465 ;
        RECT 63.510 -0.635 63.680 -0.465 ;
        RECT 65.070 -0.635 65.240 -0.465 ;
        RECT 65.430 -0.635 65.600 -0.465 ;
        RECT 65.790 -0.635 65.960 -0.465 ;
        RECT 66.150 -0.635 66.320 -0.465 ;
        RECT 66.510 -0.635 66.680 -0.465 ;
        RECT 66.870 -0.635 67.040 -0.465 ;
        RECT 68.430 -0.635 68.600 -0.465 ;
        RECT 68.790 -0.635 68.960 -0.465 ;
        RECT 69.150 -0.635 69.320 -0.465 ;
        RECT 69.510 -0.635 69.680 -0.465 ;
        RECT 69.870 -0.635 70.040 -0.465 ;
        RECT 70.230 -0.635 70.400 -0.465 ;
        RECT 71.790 -0.635 71.960 -0.465 ;
        RECT 72.150 -0.635 72.320 -0.465 ;
        RECT 72.510 -0.635 72.680 -0.465 ;
        RECT 72.870 -0.635 73.040 -0.465 ;
        RECT 73.230 -0.635 73.400 -0.465 ;
        RECT 73.590 -0.635 73.760 -0.465 ;
        RECT 75.150 -0.635 75.320 -0.465 ;
        RECT 75.510 -0.635 75.680 -0.465 ;
        RECT 75.870 -0.635 76.040 -0.465 ;
        RECT 76.230 -0.635 76.400 -0.465 ;
        RECT 76.590 -0.635 76.760 -0.465 ;
        RECT 76.950 -0.635 77.120 -0.465 ;
        RECT 78.510 -0.635 78.680 -0.465 ;
        RECT 78.870 -0.635 79.040 -0.465 ;
        RECT 79.230 -0.635 79.400 -0.465 ;
        RECT 79.590 -0.635 79.760 -0.465 ;
        RECT 79.950 -0.635 80.120 -0.465 ;
        RECT 80.310 -0.635 80.480 -0.465 ;
        RECT 81.870 -0.635 82.040 -0.465 ;
        RECT 82.230 -0.635 82.400 -0.465 ;
        RECT 82.590 -0.635 82.760 -0.465 ;
        RECT 82.950 -0.635 83.120 -0.465 ;
        RECT 83.310 -0.635 83.480 -0.465 ;
        RECT 83.670 -0.635 83.840 -0.465 ;
        RECT 85.230 -0.635 85.400 -0.465 ;
        RECT 85.590 -0.635 85.760 -0.465 ;
        RECT 85.950 -0.635 86.120 -0.465 ;
        RECT 86.310 -0.635 86.480 -0.465 ;
        RECT 86.670 -0.635 86.840 -0.465 ;
        RECT 87.030 -0.635 87.200 -0.465 ;
        RECT 88.590 -0.635 88.760 -0.465 ;
        RECT 88.950 -0.635 89.120 -0.465 ;
        RECT 89.310 -0.635 89.480 -0.465 ;
        RECT 89.670 -0.635 89.840 -0.465 ;
        RECT 90.030 -0.635 90.200 -0.465 ;
        RECT 90.390 -0.635 90.560 -0.465 ;
        RECT 91.950 -0.635 92.120 -0.465 ;
        RECT 92.310 -0.635 92.480 -0.465 ;
        RECT 92.670 -0.635 92.840 -0.465 ;
        RECT 93.030 -0.635 93.200 -0.465 ;
        RECT 93.390 -0.635 93.560 -0.465 ;
        RECT 93.750 -0.635 93.920 -0.465 ;
        RECT 95.310 -0.635 95.480 -0.465 ;
        RECT 95.670 -0.635 95.840 -0.465 ;
        RECT 96.030 -0.635 96.200 -0.465 ;
        RECT 96.390 -0.635 96.560 -0.465 ;
        RECT 96.750 -0.635 96.920 -0.465 ;
        RECT 97.110 -0.635 97.280 -0.465 ;
        RECT 98.670 -0.635 98.840 -0.465 ;
        RECT 99.030 -0.635 99.200 -0.465 ;
        RECT 99.390 -0.635 99.560 -0.465 ;
        RECT 99.750 -0.635 99.920 -0.465 ;
        RECT 100.110 -0.635 100.280 -0.465 ;
        RECT 100.470 -0.635 100.640 -0.465 ;
        RECT 102.030 -0.635 102.200 -0.465 ;
        RECT 102.390 -0.635 102.560 -0.465 ;
        RECT 102.750 -0.635 102.920 -0.465 ;
        RECT 103.110 -0.635 103.280 -0.465 ;
        RECT 103.470 -0.635 103.640 -0.465 ;
        RECT 103.830 -0.635 104.000 -0.465 ;
        RECT 105.390 -0.635 105.560 -0.465 ;
        RECT 105.750 -0.635 105.920 -0.465 ;
        RECT 106.110 -0.635 106.280 -0.465 ;
        RECT 106.470 -0.635 106.640 -0.465 ;
        RECT 106.830 -0.635 107.000 -0.465 ;
        RECT 107.190 -0.635 107.360 -0.465 ;
        RECT 108.750 -0.635 108.920 -0.465 ;
        RECT 109.110 -0.635 109.280 -0.465 ;
        RECT 109.470 -0.635 109.640 -0.465 ;
        RECT 109.830 -0.635 110.000 -0.465 ;
        RECT 110.190 -0.635 110.360 -0.465 ;
        RECT 110.550 -0.635 110.720 -0.465 ;
        RECT -2.890 -3.745 -2.720 -3.575 ;
        RECT -2.530 -3.745 -2.360 -3.575 ;
        RECT -2.170 -3.745 -2.000 -3.575 ;
        RECT -1.810 -3.745 -1.640 -3.575 ;
        RECT -1.450 -3.745 -1.280 -3.575 ;
        RECT -1.090 -3.745 -0.920 -3.575 ;
        RECT -0.730 -3.745 -0.560 -3.575 ;
        RECT 4.230 -3.745 4.400 -3.575 ;
        RECT 4.590 -3.745 4.760 -3.575 ;
        RECT 4.950 -3.745 5.120 -3.575 ;
        RECT 5.310 -3.745 5.480 -3.575 ;
        RECT 5.670 -3.745 5.840 -3.575 ;
        RECT 6.030 -3.745 6.200 -3.575 ;
        RECT 6.390 -3.745 6.560 -3.575 ;
        RECT 7.590 -3.745 7.760 -3.575 ;
        RECT 7.950 -3.745 8.120 -3.575 ;
        RECT 8.310 -3.745 8.480 -3.575 ;
        RECT 8.670 -3.745 8.840 -3.575 ;
        RECT 9.030 -3.745 9.200 -3.575 ;
        RECT 9.390 -3.745 9.560 -3.575 ;
        RECT 9.750 -3.745 9.920 -3.575 ;
        RECT 10.950 -3.745 11.120 -3.575 ;
        RECT 11.310 -3.745 11.480 -3.575 ;
        RECT 11.670 -3.745 11.840 -3.575 ;
        RECT 12.030 -3.745 12.200 -3.575 ;
        RECT 12.390 -3.745 12.560 -3.575 ;
        RECT 12.750 -3.745 12.920 -3.575 ;
        RECT 13.110 -3.745 13.280 -3.575 ;
        RECT 14.310 -3.745 14.480 -3.575 ;
        RECT 14.670 -3.745 14.840 -3.575 ;
        RECT 15.030 -3.745 15.200 -3.575 ;
        RECT 15.390 -3.745 15.560 -3.575 ;
        RECT 15.750 -3.745 15.920 -3.575 ;
        RECT 16.110 -3.745 16.280 -3.575 ;
        RECT 16.470 -3.745 16.640 -3.575 ;
        RECT 17.670 -3.745 17.840 -3.575 ;
        RECT 18.030 -3.745 18.200 -3.575 ;
        RECT 18.390 -3.745 18.560 -3.575 ;
        RECT 18.750 -3.745 18.920 -3.575 ;
        RECT 19.110 -3.745 19.280 -3.575 ;
        RECT 19.470 -3.745 19.640 -3.575 ;
        RECT 19.830 -3.745 20.000 -3.575 ;
        RECT 21.030 -3.745 21.200 -3.575 ;
        RECT 21.390 -3.745 21.560 -3.575 ;
        RECT 21.750 -3.745 21.920 -3.575 ;
        RECT 22.110 -3.745 22.280 -3.575 ;
        RECT 22.470 -3.745 22.640 -3.575 ;
        RECT 22.830 -3.745 23.000 -3.575 ;
        RECT 23.190 -3.745 23.360 -3.575 ;
        RECT 24.390 -3.745 24.560 -3.575 ;
        RECT 24.750 -3.745 24.920 -3.575 ;
        RECT 25.110 -3.745 25.280 -3.575 ;
        RECT 25.470 -3.745 25.640 -3.575 ;
        RECT 25.830 -3.745 26.000 -3.575 ;
        RECT 26.190 -3.745 26.360 -3.575 ;
        RECT 26.550 -3.745 26.720 -3.575 ;
        RECT 27.750 -3.745 27.920 -3.575 ;
        RECT 28.110 -3.745 28.280 -3.575 ;
        RECT 28.470 -3.745 28.640 -3.575 ;
        RECT 28.830 -3.745 29.000 -3.575 ;
        RECT 29.190 -3.745 29.360 -3.575 ;
        RECT 29.550 -3.745 29.720 -3.575 ;
        RECT 29.910 -3.745 30.080 -3.575 ;
        RECT 31.110 -3.745 31.280 -3.575 ;
        RECT 31.470 -3.745 31.640 -3.575 ;
        RECT 31.830 -3.745 32.000 -3.575 ;
        RECT 32.190 -3.745 32.360 -3.575 ;
        RECT 32.550 -3.745 32.720 -3.575 ;
        RECT 32.910 -3.745 33.080 -3.575 ;
        RECT 33.270 -3.745 33.440 -3.575 ;
        RECT 34.470 -3.745 34.640 -3.575 ;
        RECT 34.830 -3.745 35.000 -3.575 ;
        RECT 35.190 -3.745 35.360 -3.575 ;
        RECT 35.550 -3.745 35.720 -3.575 ;
        RECT 35.910 -3.745 36.080 -3.575 ;
        RECT 36.270 -3.745 36.440 -3.575 ;
        RECT 36.630 -3.745 36.800 -3.575 ;
        RECT 37.830 -3.745 38.000 -3.575 ;
        RECT 38.190 -3.745 38.360 -3.575 ;
        RECT 38.550 -3.745 38.720 -3.575 ;
        RECT 38.910 -3.745 39.080 -3.575 ;
        RECT 39.270 -3.745 39.440 -3.575 ;
        RECT 39.630 -3.745 39.800 -3.575 ;
        RECT 39.990 -3.745 40.160 -3.575 ;
        RECT 41.190 -3.745 41.360 -3.575 ;
        RECT 41.550 -3.745 41.720 -3.575 ;
        RECT 41.910 -3.745 42.080 -3.575 ;
        RECT 42.270 -3.745 42.440 -3.575 ;
        RECT 42.630 -3.745 42.800 -3.575 ;
        RECT 42.990 -3.745 43.160 -3.575 ;
        RECT 43.350 -3.745 43.520 -3.575 ;
        RECT 44.550 -3.745 44.720 -3.575 ;
        RECT 44.910 -3.745 45.080 -3.575 ;
        RECT 45.270 -3.745 45.440 -3.575 ;
        RECT 45.630 -3.745 45.800 -3.575 ;
        RECT 45.990 -3.745 46.160 -3.575 ;
        RECT 46.350 -3.745 46.520 -3.575 ;
        RECT 46.710 -3.745 46.880 -3.575 ;
        RECT 47.910 -3.745 48.080 -3.575 ;
        RECT 48.270 -3.745 48.440 -3.575 ;
        RECT 48.630 -3.745 48.800 -3.575 ;
        RECT 48.990 -3.745 49.160 -3.575 ;
        RECT 49.350 -3.745 49.520 -3.575 ;
        RECT 49.710 -3.745 49.880 -3.575 ;
        RECT 50.070 -3.745 50.240 -3.575 ;
        RECT 51.270 -3.745 51.440 -3.575 ;
        RECT 51.630 -3.745 51.800 -3.575 ;
        RECT 51.990 -3.745 52.160 -3.575 ;
        RECT 52.350 -3.745 52.520 -3.575 ;
        RECT 52.710 -3.745 52.880 -3.575 ;
        RECT 53.070 -3.745 53.240 -3.575 ;
        RECT 53.430 -3.745 53.600 -3.575 ;
        RECT 54.630 -3.745 54.800 -3.575 ;
        RECT 54.990 -3.745 55.160 -3.575 ;
        RECT 55.350 -3.745 55.520 -3.575 ;
        RECT 55.710 -3.745 55.880 -3.575 ;
        RECT 56.070 -3.745 56.240 -3.575 ;
        RECT 56.430 -3.745 56.600 -3.575 ;
        RECT 56.790 -3.745 56.960 -3.575 ;
        RECT 57.990 -3.745 58.160 -3.575 ;
        RECT 58.350 -3.745 58.520 -3.575 ;
        RECT 58.710 -3.745 58.880 -3.575 ;
        RECT 59.070 -3.745 59.240 -3.575 ;
        RECT 59.430 -3.745 59.600 -3.575 ;
        RECT 59.790 -3.745 59.960 -3.575 ;
        RECT 60.150 -3.745 60.320 -3.575 ;
        RECT 61.350 -3.745 61.520 -3.575 ;
        RECT 61.710 -3.745 61.880 -3.575 ;
        RECT 62.070 -3.745 62.240 -3.575 ;
        RECT 62.430 -3.745 62.600 -3.575 ;
        RECT 62.790 -3.745 62.960 -3.575 ;
        RECT 63.150 -3.745 63.320 -3.575 ;
        RECT 63.510 -3.745 63.680 -3.575 ;
        RECT 64.710 -3.745 64.880 -3.575 ;
        RECT 65.070 -3.745 65.240 -3.575 ;
        RECT 65.430 -3.745 65.600 -3.575 ;
        RECT 65.790 -3.745 65.960 -3.575 ;
        RECT 66.150 -3.745 66.320 -3.575 ;
        RECT 66.510 -3.745 66.680 -3.575 ;
        RECT 66.870 -3.745 67.040 -3.575 ;
        RECT 68.070 -3.745 68.240 -3.575 ;
        RECT 68.430 -3.745 68.600 -3.575 ;
        RECT 68.790 -3.745 68.960 -3.575 ;
        RECT 69.150 -3.745 69.320 -3.575 ;
        RECT 69.510 -3.745 69.680 -3.575 ;
        RECT 69.870 -3.745 70.040 -3.575 ;
        RECT 70.230 -3.745 70.400 -3.575 ;
        RECT 71.430 -3.745 71.600 -3.575 ;
        RECT 71.790 -3.745 71.960 -3.575 ;
        RECT 72.150 -3.745 72.320 -3.575 ;
        RECT 72.510 -3.745 72.680 -3.575 ;
        RECT 72.870 -3.745 73.040 -3.575 ;
        RECT 73.230 -3.745 73.400 -3.575 ;
        RECT 73.590 -3.745 73.760 -3.575 ;
        RECT 74.790 -3.745 74.960 -3.575 ;
        RECT 75.150 -3.745 75.320 -3.575 ;
        RECT 75.510 -3.745 75.680 -3.575 ;
        RECT 75.870 -3.745 76.040 -3.575 ;
        RECT 76.230 -3.745 76.400 -3.575 ;
        RECT 76.590 -3.745 76.760 -3.575 ;
        RECT 76.950 -3.745 77.120 -3.575 ;
        RECT 78.150 -3.745 78.320 -3.575 ;
        RECT 78.510 -3.745 78.680 -3.575 ;
        RECT 78.870 -3.745 79.040 -3.575 ;
        RECT 79.230 -3.745 79.400 -3.575 ;
        RECT 79.590 -3.745 79.760 -3.575 ;
        RECT 79.950 -3.745 80.120 -3.575 ;
        RECT 80.310 -3.745 80.480 -3.575 ;
        RECT 81.510 -3.745 81.680 -3.575 ;
        RECT 81.870 -3.745 82.040 -3.575 ;
        RECT 82.230 -3.745 82.400 -3.575 ;
        RECT 82.590 -3.745 82.760 -3.575 ;
        RECT 82.950 -3.745 83.120 -3.575 ;
        RECT 83.310 -3.745 83.480 -3.575 ;
        RECT 83.670 -3.745 83.840 -3.575 ;
        RECT 84.870 -3.745 85.040 -3.575 ;
        RECT 85.230 -3.745 85.400 -3.575 ;
        RECT 85.590 -3.745 85.760 -3.575 ;
        RECT 85.950 -3.745 86.120 -3.575 ;
        RECT 86.310 -3.745 86.480 -3.575 ;
        RECT 86.670 -3.745 86.840 -3.575 ;
        RECT 87.030 -3.745 87.200 -3.575 ;
        RECT 88.230 -3.745 88.400 -3.575 ;
        RECT 88.590 -3.745 88.760 -3.575 ;
        RECT 88.950 -3.745 89.120 -3.575 ;
        RECT 89.310 -3.745 89.480 -3.575 ;
        RECT 89.670 -3.745 89.840 -3.575 ;
        RECT 90.030 -3.745 90.200 -3.575 ;
        RECT 90.390 -3.745 90.560 -3.575 ;
        RECT 91.590 -3.745 91.760 -3.575 ;
        RECT 91.950 -3.745 92.120 -3.575 ;
        RECT 92.310 -3.745 92.480 -3.575 ;
        RECT 92.670 -3.745 92.840 -3.575 ;
        RECT 93.030 -3.745 93.200 -3.575 ;
        RECT 93.390 -3.745 93.560 -3.575 ;
        RECT 93.750 -3.745 93.920 -3.575 ;
        RECT 94.950 -3.745 95.120 -3.575 ;
        RECT 95.310 -3.745 95.480 -3.575 ;
        RECT 95.670 -3.745 95.840 -3.575 ;
        RECT 96.030 -3.745 96.200 -3.575 ;
        RECT 96.390 -3.745 96.560 -3.575 ;
        RECT 96.750 -3.745 96.920 -3.575 ;
        RECT 97.110 -3.745 97.280 -3.575 ;
        RECT 98.310 -3.745 98.480 -3.575 ;
        RECT 98.670 -3.745 98.840 -3.575 ;
        RECT 99.030 -3.745 99.200 -3.575 ;
        RECT 99.390 -3.745 99.560 -3.575 ;
        RECT 99.750 -3.745 99.920 -3.575 ;
        RECT 100.110 -3.745 100.280 -3.575 ;
        RECT 100.470 -3.745 100.640 -3.575 ;
        RECT 101.670 -3.745 101.840 -3.575 ;
        RECT 102.030 -3.745 102.200 -3.575 ;
        RECT 102.390 -3.745 102.560 -3.575 ;
        RECT 102.750 -3.745 102.920 -3.575 ;
        RECT 103.110 -3.745 103.280 -3.575 ;
        RECT 103.470 -3.745 103.640 -3.575 ;
        RECT 103.830 -3.745 104.000 -3.575 ;
        RECT 105.030 -3.745 105.200 -3.575 ;
        RECT 105.390 -3.745 105.560 -3.575 ;
        RECT 105.750 -3.745 105.920 -3.575 ;
        RECT 106.110 -3.745 106.280 -3.575 ;
        RECT 106.470 -3.745 106.640 -3.575 ;
        RECT 106.830 -3.745 107.000 -3.575 ;
        RECT 107.190 -3.745 107.360 -3.575 ;
        RECT 108.390 -3.745 108.560 -3.575 ;
        RECT 108.750 -3.745 108.920 -3.575 ;
        RECT 109.110 -3.745 109.280 -3.575 ;
        RECT 109.470 -3.745 109.640 -3.575 ;
        RECT 109.830 -3.745 110.000 -3.575 ;
        RECT 110.190 -3.745 110.360 -3.575 ;
        RECT 110.550 -3.745 110.720 -3.575 ;
        RECT -3.205 -4.225 -3.035 -4.055 ;
        RECT -2.725 -4.225 -2.555 -4.055 ;
        RECT -2.245 -4.225 -2.075 -4.055 ;
        RECT -1.765 -4.225 -1.595 -4.055 ;
        RECT -1.285 -4.225 -1.115 -4.055 ;
        RECT -0.805 -4.225 -0.635 -4.055 ;
        RECT -0.325 -4.225 -0.155 -4.055 ;
        RECT 3.915 -4.225 4.085 -4.055 ;
        RECT 4.395 -4.225 4.565 -4.055 ;
        RECT 4.875 -4.225 5.045 -4.055 ;
        RECT 5.355 -4.225 5.525 -4.055 ;
        RECT 5.835 -4.225 6.005 -4.055 ;
        RECT 6.315 -4.225 6.485 -4.055 ;
        RECT 6.795 -4.225 6.965 -4.055 ;
        RECT 7.275 -4.225 7.445 -4.055 ;
        RECT 7.755 -4.225 7.925 -4.055 ;
        RECT 8.235 -4.225 8.405 -4.055 ;
        RECT 8.715 -4.225 8.885 -4.055 ;
        RECT 9.195 -4.225 9.365 -4.055 ;
        RECT 9.675 -4.225 9.845 -4.055 ;
        RECT 10.155 -4.225 10.325 -4.055 ;
        RECT 10.635 -4.225 10.805 -4.055 ;
        RECT 11.115 -4.225 11.285 -4.055 ;
        RECT 11.595 -4.225 11.765 -4.055 ;
        RECT 12.075 -4.225 12.245 -4.055 ;
        RECT 12.555 -4.225 12.725 -4.055 ;
        RECT 13.035 -4.225 13.205 -4.055 ;
        RECT 13.515 -4.225 13.685 -4.055 ;
        RECT 13.995 -4.225 14.165 -4.055 ;
        RECT 14.475 -4.225 14.645 -4.055 ;
        RECT 14.955 -4.225 15.125 -4.055 ;
        RECT 15.435 -4.225 15.605 -4.055 ;
        RECT 15.915 -4.225 16.085 -4.055 ;
        RECT 16.395 -4.225 16.565 -4.055 ;
        RECT 16.875 -4.225 17.045 -4.055 ;
        RECT 17.355 -4.225 17.525 -4.055 ;
        RECT 17.835 -4.225 18.005 -4.055 ;
        RECT 18.315 -4.225 18.485 -4.055 ;
        RECT 18.795 -4.225 18.965 -4.055 ;
        RECT 19.275 -4.225 19.445 -4.055 ;
        RECT 19.755 -4.225 19.925 -4.055 ;
        RECT 20.235 -4.225 20.405 -4.055 ;
        RECT 20.715 -4.225 20.885 -4.055 ;
        RECT 21.195 -4.225 21.365 -4.055 ;
        RECT 21.675 -4.225 21.845 -4.055 ;
        RECT 22.155 -4.225 22.325 -4.055 ;
        RECT 22.635 -4.225 22.805 -4.055 ;
        RECT 23.115 -4.225 23.285 -4.055 ;
        RECT 23.595 -4.225 23.765 -4.055 ;
        RECT 24.075 -4.225 24.245 -4.055 ;
        RECT 24.555 -4.225 24.725 -4.055 ;
        RECT 25.035 -4.225 25.205 -4.055 ;
        RECT 25.515 -4.225 25.685 -4.055 ;
        RECT 25.995 -4.225 26.165 -4.055 ;
        RECT 26.475 -4.225 26.645 -4.055 ;
        RECT 26.955 -4.225 27.125 -4.055 ;
        RECT 27.435 -4.225 27.605 -4.055 ;
        RECT 27.915 -4.225 28.085 -4.055 ;
        RECT 28.395 -4.225 28.565 -4.055 ;
        RECT 28.875 -4.225 29.045 -4.055 ;
        RECT 29.355 -4.225 29.525 -4.055 ;
        RECT 29.835 -4.225 30.005 -4.055 ;
        RECT 30.315 -4.225 30.485 -4.055 ;
        RECT 30.795 -4.225 30.965 -4.055 ;
        RECT 31.275 -4.225 31.445 -4.055 ;
        RECT 31.755 -4.225 31.925 -4.055 ;
        RECT 32.235 -4.225 32.405 -4.055 ;
        RECT 32.715 -4.225 32.885 -4.055 ;
        RECT 33.195 -4.225 33.365 -4.055 ;
        RECT 33.675 -4.225 33.845 -4.055 ;
        RECT 34.155 -4.225 34.325 -4.055 ;
        RECT 34.635 -4.225 34.805 -4.055 ;
        RECT 35.115 -4.225 35.285 -4.055 ;
        RECT 35.595 -4.225 35.765 -4.055 ;
        RECT 36.075 -4.225 36.245 -4.055 ;
        RECT 36.555 -4.225 36.725 -4.055 ;
        RECT 37.035 -4.225 37.205 -4.055 ;
        RECT 37.515 -4.225 37.685 -4.055 ;
        RECT 37.995 -4.225 38.165 -4.055 ;
        RECT 38.475 -4.225 38.645 -4.055 ;
        RECT 38.955 -4.225 39.125 -4.055 ;
        RECT 39.435 -4.225 39.605 -4.055 ;
        RECT 39.915 -4.225 40.085 -4.055 ;
        RECT 40.395 -4.225 40.565 -4.055 ;
        RECT 40.875 -4.225 41.045 -4.055 ;
        RECT 41.355 -4.225 41.525 -4.055 ;
        RECT 41.835 -4.225 42.005 -4.055 ;
        RECT 42.315 -4.225 42.485 -4.055 ;
        RECT 42.795 -4.225 42.965 -4.055 ;
        RECT 43.275 -4.225 43.445 -4.055 ;
        RECT 43.755 -4.225 43.925 -4.055 ;
        RECT 44.235 -4.225 44.405 -4.055 ;
        RECT 44.715 -4.225 44.885 -4.055 ;
        RECT 45.195 -4.225 45.365 -4.055 ;
        RECT 45.675 -4.225 45.845 -4.055 ;
        RECT 46.155 -4.225 46.325 -4.055 ;
        RECT 46.635 -4.225 46.805 -4.055 ;
        RECT 47.115 -4.225 47.285 -4.055 ;
        RECT 47.595 -4.225 47.765 -4.055 ;
        RECT 48.075 -4.225 48.245 -4.055 ;
        RECT 48.555 -4.225 48.725 -4.055 ;
        RECT 49.035 -4.225 49.205 -4.055 ;
        RECT 49.515 -4.225 49.685 -4.055 ;
        RECT 49.995 -4.225 50.165 -4.055 ;
        RECT 50.475 -4.225 50.645 -4.055 ;
        RECT 50.955 -4.225 51.125 -4.055 ;
        RECT 51.435 -4.225 51.605 -4.055 ;
        RECT 51.915 -4.225 52.085 -4.055 ;
        RECT 52.395 -4.225 52.565 -4.055 ;
        RECT 52.875 -4.225 53.045 -4.055 ;
        RECT 53.355 -4.225 53.525 -4.055 ;
        RECT 53.835 -4.225 54.005 -4.055 ;
        RECT 54.315 -4.225 54.485 -4.055 ;
        RECT 54.795 -4.225 54.965 -4.055 ;
        RECT 55.275 -4.225 55.445 -4.055 ;
        RECT 55.755 -4.225 55.925 -4.055 ;
        RECT 56.235 -4.225 56.405 -4.055 ;
        RECT 56.715 -4.225 56.885 -4.055 ;
        RECT 57.195 -4.225 57.365 -4.055 ;
        RECT 57.675 -4.225 57.845 -4.055 ;
        RECT 58.155 -4.225 58.325 -4.055 ;
        RECT 58.635 -4.225 58.805 -4.055 ;
        RECT 59.115 -4.225 59.285 -4.055 ;
        RECT 59.595 -4.225 59.765 -4.055 ;
        RECT 60.075 -4.225 60.245 -4.055 ;
        RECT 60.555 -4.225 60.725 -4.055 ;
        RECT 61.035 -4.225 61.205 -4.055 ;
        RECT 61.515 -4.225 61.685 -4.055 ;
        RECT 61.995 -4.225 62.165 -4.055 ;
        RECT 62.475 -4.225 62.645 -4.055 ;
        RECT 62.955 -4.225 63.125 -4.055 ;
        RECT 63.435 -4.225 63.605 -4.055 ;
        RECT 63.915 -4.225 64.085 -4.055 ;
        RECT 64.395 -4.225 64.565 -4.055 ;
        RECT 64.875 -4.225 65.045 -4.055 ;
        RECT 65.355 -4.225 65.525 -4.055 ;
        RECT 65.835 -4.225 66.005 -4.055 ;
        RECT 66.315 -4.225 66.485 -4.055 ;
        RECT 66.795 -4.225 66.965 -4.055 ;
        RECT 67.275 -4.225 67.445 -4.055 ;
        RECT 67.755 -4.225 67.925 -4.055 ;
        RECT 68.235 -4.225 68.405 -4.055 ;
        RECT 68.715 -4.225 68.885 -4.055 ;
        RECT 69.195 -4.225 69.365 -4.055 ;
        RECT 69.675 -4.225 69.845 -4.055 ;
        RECT 70.155 -4.225 70.325 -4.055 ;
        RECT 70.635 -4.225 70.805 -4.055 ;
        RECT 71.115 -4.225 71.285 -4.055 ;
        RECT 71.595 -4.225 71.765 -4.055 ;
        RECT 72.075 -4.225 72.245 -4.055 ;
        RECT 72.555 -4.225 72.725 -4.055 ;
        RECT 73.035 -4.225 73.205 -4.055 ;
        RECT 73.515 -4.225 73.685 -4.055 ;
        RECT 73.995 -4.225 74.165 -4.055 ;
        RECT 74.475 -4.225 74.645 -4.055 ;
        RECT 74.955 -4.225 75.125 -4.055 ;
        RECT 75.435 -4.225 75.605 -4.055 ;
        RECT 75.915 -4.225 76.085 -4.055 ;
        RECT 76.395 -4.225 76.565 -4.055 ;
        RECT 76.875 -4.225 77.045 -4.055 ;
        RECT 77.355 -4.225 77.525 -4.055 ;
        RECT 77.835 -4.225 78.005 -4.055 ;
        RECT 78.315 -4.225 78.485 -4.055 ;
        RECT 78.795 -4.225 78.965 -4.055 ;
        RECT 79.275 -4.225 79.445 -4.055 ;
        RECT 79.755 -4.225 79.925 -4.055 ;
        RECT 80.235 -4.225 80.405 -4.055 ;
        RECT 80.715 -4.225 80.885 -4.055 ;
        RECT 81.195 -4.225 81.365 -4.055 ;
        RECT 81.675 -4.225 81.845 -4.055 ;
        RECT 82.155 -4.225 82.325 -4.055 ;
        RECT 82.635 -4.225 82.805 -4.055 ;
        RECT 83.115 -4.225 83.285 -4.055 ;
        RECT 83.595 -4.225 83.765 -4.055 ;
        RECT 84.075 -4.225 84.245 -4.055 ;
        RECT 84.555 -4.225 84.725 -4.055 ;
        RECT 85.035 -4.225 85.205 -4.055 ;
        RECT 85.515 -4.225 85.685 -4.055 ;
        RECT 85.995 -4.225 86.165 -4.055 ;
        RECT 86.475 -4.225 86.645 -4.055 ;
        RECT 86.955 -4.225 87.125 -4.055 ;
        RECT 87.435 -4.225 87.605 -4.055 ;
        RECT 87.915 -4.225 88.085 -4.055 ;
        RECT 88.395 -4.225 88.565 -4.055 ;
        RECT 88.875 -4.225 89.045 -4.055 ;
        RECT 89.355 -4.225 89.525 -4.055 ;
        RECT 89.835 -4.225 90.005 -4.055 ;
        RECT 90.315 -4.225 90.485 -4.055 ;
        RECT 90.795 -4.225 90.965 -4.055 ;
        RECT 91.275 -4.225 91.445 -4.055 ;
        RECT 91.755 -4.225 91.925 -4.055 ;
        RECT 92.235 -4.225 92.405 -4.055 ;
        RECT 92.715 -4.225 92.885 -4.055 ;
        RECT 93.195 -4.225 93.365 -4.055 ;
        RECT 93.675 -4.225 93.845 -4.055 ;
        RECT 94.155 -4.225 94.325 -4.055 ;
        RECT 94.635 -4.225 94.805 -4.055 ;
        RECT 95.115 -4.225 95.285 -4.055 ;
        RECT 95.595 -4.225 95.765 -4.055 ;
        RECT 96.075 -4.225 96.245 -4.055 ;
        RECT 96.555 -4.225 96.725 -4.055 ;
        RECT 97.035 -4.225 97.205 -4.055 ;
        RECT 97.515 -4.225 97.685 -4.055 ;
        RECT 97.995 -4.225 98.165 -4.055 ;
        RECT 98.475 -4.225 98.645 -4.055 ;
        RECT 98.955 -4.225 99.125 -4.055 ;
        RECT 99.435 -4.225 99.605 -4.055 ;
        RECT 99.915 -4.225 100.085 -4.055 ;
        RECT 100.395 -4.225 100.565 -4.055 ;
        RECT 100.875 -4.225 101.045 -4.055 ;
        RECT 101.355 -4.225 101.525 -4.055 ;
        RECT 101.835 -4.225 102.005 -4.055 ;
        RECT 102.315 -4.225 102.485 -4.055 ;
        RECT 102.795 -4.225 102.965 -4.055 ;
        RECT 103.275 -4.225 103.445 -4.055 ;
        RECT 103.755 -4.225 103.925 -4.055 ;
        RECT 104.235 -4.225 104.405 -4.055 ;
        RECT 104.715 -4.225 104.885 -4.055 ;
        RECT 105.195 -4.225 105.365 -4.055 ;
        RECT 105.675 -4.225 105.845 -4.055 ;
        RECT 106.155 -4.225 106.325 -4.055 ;
        RECT 106.635 -4.225 106.805 -4.055 ;
        RECT 107.115 -4.225 107.285 -4.055 ;
        RECT 107.595 -4.225 107.765 -4.055 ;
        RECT 108.075 -4.225 108.245 -4.055 ;
        RECT 108.555 -4.225 108.725 -4.055 ;
        RECT 109.035 -4.225 109.205 -4.055 ;
        RECT 109.515 -4.225 109.685 -4.055 ;
        RECT 109.995 -4.225 110.165 -4.055 ;
        RECT 110.475 -4.225 110.645 -4.055 ;
        RECT 110.955 -4.225 111.125 -4.055 ;
      LAYER met1 ;
        RECT -3.360 3.375 0.000 4.120 ;
        RECT 2.030 -0.690 111.280 0.050 ;
        RECT 3.760 -0.695 111.280 -0.690 ;
        RECT -3.360 -3.630 0.000 -3.515 ;
        RECT 3.760 -3.630 111.280 -3.515 ;
        RECT -3.360 -4.170 111.280 -3.630 ;
        RECT -3.360 -4.255 0.000 -4.170 ;
        RECT 3.760 -4.255 111.280 -4.170 ;
  END
END wl_driver
END LIBRARY

